
module global_buffer_0 ( clk, rst, wr_en, index, data_in, data_out );
  input [7:0] index;
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, wr_en;
  wire   N10, N11, N12, N13, N14, \gbuff[1][31] , \gbuff[1][30] ,
         \gbuff[1][29] , \gbuff[1][28] , \gbuff[1][27] , \gbuff[1][26] ,
         \gbuff[1][25] , \gbuff[1][24] , \gbuff[1][23] , \gbuff[1][22] ,
         \gbuff[1][21] , \gbuff[1][20] , \gbuff[1][19] , \gbuff[1][18] ,
         \gbuff[1][17] , \gbuff[1][16] , \gbuff[1][15] , \gbuff[1][14] ,
         \gbuff[1][13] , \gbuff[1][12] , \gbuff[1][11] , \gbuff[1][10] ,
         \gbuff[1][9] , \gbuff[1][8] , \gbuff[1][7] , \gbuff[1][6] ,
         \gbuff[1][5] , \gbuff[1][4] , \gbuff[1][3] , \gbuff[1][2] ,
         \gbuff[1][1] , \gbuff[1][0] , \gbuff[0][31] , \gbuff[0][30] ,
         \gbuff[0][29] , \gbuff[0][28] , \gbuff[0][27] , \gbuff[0][26] ,
         \gbuff[0][25] , \gbuff[0][24] , \gbuff[0][23] , \gbuff[0][22] ,
         \gbuff[0][21] , \gbuff[0][20] , \gbuff[0][19] , \gbuff[0][18] ,
         \gbuff[0][17] , \gbuff[0][16] , \gbuff[0][15] , \gbuff[0][14] ,
         \gbuff[0][13] , \gbuff[0][12] , \gbuff[0][11] , \gbuff[0][10] ,
         \gbuff[0][9] , \gbuff[0][8] , \gbuff[0][7] , \gbuff[0][6] ,
         \gbuff[0][5] , \gbuff[0][4] , \gbuff[0][3] , \gbuff[0][2] ,
         \gbuff[0][1] , \gbuff[0][0] , \gbuff[3][31] , \gbuff[3][30] ,
         \gbuff[3][29] , \gbuff[3][28] , \gbuff[3][27] , \gbuff[3][26] ,
         \gbuff[3][25] , \gbuff[3][24] , \gbuff[3][23] , \gbuff[3][22] ,
         \gbuff[3][21] , \gbuff[3][20] , \gbuff[3][19] , \gbuff[3][18] ,
         \gbuff[3][17] , \gbuff[3][16] , \gbuff[3][15] , \gbuff[3][14] ,
         \gbuff[3][13] , \gbuff[3][12] , \gbuff[3][11] , \gbuff[3][10] ,
         \gbuff[3][9] , \gbuff[3][8] , \gbuff[3][7] , \gbuff[3][6] ,
         \gbuff[3][5] , \gbuff[3][4] , \gbuff[3][3] , \gbuff[3][2] ,
         \gbuff[3][1] , \gbuff[3][0] , \gbuff[2][31] , \gbuff[2][30] ,
         \gbuff[2][29] , \gbuff[2][28] , \gbuff[2][27] , \gbuff[2][26] ,
         \gbuff[2][25] , \gbuff[2][24] , \gbuff[2][23] , \gbuff[2][22] ,
         \gbuff[2][21] , \gbuff[2][20] , \gbuff[2][19] , \gbuff[2][18] ,
         \gbuff[2][17] , \gbuff[2][16] , \gbuff[2][15] , \gbuff[2][14] ,
         \gbuff[2][13] , \gbuff[2][12] , \gbuff[2][11] , \gbuff[2][10] ,
         \gbuff[2][9] , \gbuff[2][8] , \gbuff[2][7] , \gbuff[2][6] ,
         \gbuff[2][5] , \gbuff[2][4] , \gbuff[2][3] , \gbuff[2][2] ,
         \gbuff[2][1] , \gbuff[2][0] , \gbuff[5][31] , \gbuff[5][30] ,
         \gbuff[5][29] , \gbuff[5][28] , \gbuff[5][27] , \gbuff[5][26] ,
         \gbuff[5][25] , \gbuff[5][24] , \gbuff[5][23] , \gbuff[5][22] ,
         \gbuff[5][21] , \gbuff[5][20] , \gbuff[5][19] , \gbuff[5][18] ,
         \gbuff[5][17] , \gbuff[5][16] , \gbuff[5][15] , \gbuff[5][14] ,
         \gbuff[5][13] , \gbuff[5][12] , \gbuff[5][11] , \gbuff[5][10] ,
         \gbuff[5][9] , \gbuff[5][8] , \gbuff[5][7] , \gbuff[5][6] ,
         \gbuff[5][5] , \gbuff[5][4] , \gbuff[5][3] , \gbuff[5][2] ,
         \gbuff[5][1] , \gbuff[5][0] , \gbuff[4][31] , \gbuff[4][30] ,
         \gbuff[4][29] , \gbuff[4][28] , \gbuff[4][27] , \gbuff[4][26] ,
         \gbuff[4][25] , \gbuff[4][24] , \gbuff[4][23] , \gbuff[4][22] ,
         \gbuff[4][21] , \gbuff[4][20] , \gbuff[4][19] , \gbuff[4][18] ,
         \gbuff[4][17] , \gbuff[4][16] , \gbuff[4][15] , \gbuff[4][14] ,
         \gbuff[4][13] , \gbuff[4][12] , \gbuff[4][11] , \gbuff[4][10] ,
         \gbuff[4][9] , \gbuff[4][8] , \gbuff[4][7] , \gbuff[4][6] ,
         \gbuff[4][5] , \gbuff[4][4] , \gbuff[4][3] , \gbuff[4][2] ,
         \gbuff[4][1] , \gbuff[4][0] , \gbuff[7][31] , \gbuff[7][30] ,
         \gbuff[7][29] , \gbuff[7][28] , \gbuff[7][27] , \gbuff[7][26] ,
         \gbuff[7][25] , \gbuff[7][24] , \gbuff[7][23] , \gbuff[7][22] ,
         \gbuff[7][21] , \gbuff[7][20] , \gbuff[7][19] , \gbuff[7][18] ,
         \gbuff[7][17] , \gbuff[7][16] , \gbuff[7][15] , \gbuff[7][14] ,
         \gbuff[7][13] , \gbuff[7][12] , \gbuff[7][11] , \gbuff[7][10] ,
         \gbuff[7][9] , \gbuff[7][8] , \gbuff[7][7] , \gbuff[7][6] ,
         \gbuff[7][5] , \gbuff[7][4] , \gbuff[7][3] , \gbuff[7][2] ,
         \gbuff[7][1] , \gbuff[7][0] , \gbuff[6][31] , \gbuff[6][30] ,
         \gbuff[6][29] , \gbuff[6][28] , \gbuff[6][27] , \gbuff[6][26] ,
         \gbuff[6][25] , \gbuff[6][24] , \gbuff[6][23] , \gbuff[6][22] ,
         \gbuff[6][21] , \gbuff[6][20] , \gbuff[6][19] , \gbuff[6][18] ,
         \gbuff[6][17] , \gbuff[6][16] , \gbuff[6][15] , \gbuff[6][14] ,
         \gbuff[6][13] , \gbuff[6][12] , \gbuff[6][11] , \gbuff[6][10] ,
         \gbuff[6][9] , \gbuff[6][8] , \gbuff[6][7] , \gbuff[6][6] ,
         \gbuff[6][5] , \gbuff[6][4] , \gbuff[6][3] , \gbuff[6][2] ,
         \gbuff[6][1] , \gbuff[6][0] , \gbuff[9][31] , \gbuff[9][30] ,
         \gbuff[9][29] , \gbuff[9][28] , \gbuff[9][27] , \gbuff[9][26] ,
         \gbuff[9][25] , \gbuff[9][24] , \gbuff[9][23] , \gbuff[9][22] ,
         \gbuff[9][21] , \gbuff[9][20] , \gbuff[9][19] , \gbuff[9][18] ,
         \gbuff[9][17] , \gbuff[9][16] , \gbuff[9][15] , \gbuff[9][14] ,
         \gbuff[9][13] , \gbuff[9][12] , \gbuff[9][11] , \gbuff[9][10] ,
         \gbuff[9][9] , \gbuff[9][8] , \gbuff[9][7] , \gbuff[9][6] ,
         \gbuff[9][5] , \gbuff[9][4] , \gbuff[9][3] , \gbuff[9][2] ,
         \gbuff[9][1] , \gbuff[9][0] , \gbuff[8][31] , \gbuff[8][30] ,
         \gbuff[8][29] , \gbuff[8][28] , \gbuff[8][27] , \gbuff[8][26] ,
         \gbuff[8][25] , \gbuff[8][24] , \gbuff[8][23] , \gbuff[8][22] ,
         \gbuff[8][21] , \gbuff[8][20] , \gbuff[8][19] , \gbuff[8][18] ,
         \gbuff[8][17] , \gbuff[8][16] , \gbuff[8][15] , \gbuff[8][14] ,
         \gbuff[8][13] , \gbuff[8][12] , \gbuff[8][11] , \gbuff[8][10] ,
         \gbuff[8][9] , \gbuff[8][8] , \gbuff[8][7] , \gbuff[8][6] ,
         \gbuff[8][5] , \gbuff[8][4] , \gbuff[8][3] , \gbuff[8][2] ,
         \gbuff[8][1] , \gbuff[8][0] , \gbuff[11][31] , \gbuff[11][30] ,
         \gbuff[11][29] , \gbuff[11][28] , \gbuff[11][27] , \gbuff[11][26] ,
         \gbuff[11][25] , \gbuff[11][24] , \gbuff[11][23] , \gbuff[11][22] ,
         \gbuff[11][21] , \gbuff[11][20] , \gbuff[11][19] , \gbuff[11][18] ,
         \gbuff[11][17] , \gbuff[11][16] , \gbuff[11][15] , \gbuff[11][14] ,
         \gbuff[11][13] , \gbuff[11][12] , \gbuff[11][11] , \gbuff[11][10] ,
         \gbuff[11][9] , \gbuff[11][8] , \gbuff[11][7] , \gbuff[11][6] ,
         \gbuff[11][5] , \gbuff[11][4] , \gbuff[11][3] , \gbuff[11][2] ,
         \gbuff[11][1] , \gbuff[11][0] , \gbuff[10][31] , \gbuff[10][30] ,
         \gbuff[10][29] , \gbuff[10][28] , \gbuff[10][27] , \gbuff[10][26] ,
         \gbuff[10][25] , \gbuff[10][24] , \gbuff[10][23] , \gbuff[10][22] ,
         \gbuff[10][21] , \gbuff[10][20] , \gbuff[10][19] , \gbuff[10][18] ,
         \gbuff[10][17] , \gbuff[10][16] , \gbuff[10][15] , \gbuff[10][14] ,
         \gbuff[10][13] , \gbuff[10][12] , \gbuff[10][11] , \gbuff[10][10] ,
         \gbuff[10][9] , \gbuff[10][8] , \gbuff[10][7] , \gbuff[10][6] ,
         \gbuff[10][5] , \gbuff[10][4] , \gbuff[10][3] , \gbuff[10][2] ,
         \gbuff[10][1] , \gbuff[10][0] , \gbuff[13][31] , \gbuff[13][30] ,
         \gbuff[13][29] , \gbuff[13][28] , \gbuff[13][27] , \gbuff[13][26] ,
         \gbuff[13][25] , \gbuff[13][24] , \gbuff[13][23] , \gbuff[13][22] ,
         \gbuff[13][21] , \gbuff[13][20] , \gbuff[13][19] , \gbuff[13][18] ,
         \gbuff[13][17] , \gbuff[13][16] , \gbuff[13][15] , \gbuff[13][14] ,
         \gbuff[13][13] , \gbuff[13][12] , \gbuff[13][11] , \gbuff[13][10] ,
         \gbuff[13][9] , \gbuff[13][8] , \gbuff[13][7] , \gbuff[13][6] ,
         \gbuff[13][5] , \gbuff[13][4] , \gbuff[13][3] , \gbuff[13][2] ,
         \gbuff[13][1] , \gbuff[13][0] , \gbuff[12][31] , \gbuff[12][30] ,
         \gbuff[12][29] , \gbuff[12][28] , \gbuff[12][27] , \gbuff[12][26] ,
         \gbuff[12][25] , \gbuff[12][24] , \gbuff[12][23] , \gbuff[12][22] ,
         \gbuff[12][21] , \gbuff[12][20] , \gbuff[12][19] , \gbuff[12][18] ,
         \gbuff[12][17] , \gbuff[12][16] , \gbuff[12][15] , \gbuff[12][14] ,
         \gbuff[12][13] , \gbuff[12][12] , \gbuff[12][11] , \gbuff[12][10] ,
         \gbuff[12][9] , \gbuff[12][8] , \gbuff[12][7] , \gbuff[12][6] ,
         \gbuff[12][5] , \gbuff[12][4] , \gbuff[12][3] , \gbuff[12][2] ,
         \gbuff[12][1] , \gbuff[12][0] , \gbuff[15][31] , \gbuff[15][30] ,
         \gbuff[15][29] , \gbuff[15][28] , \gbuff[15][27] , \gbuff[15][26] ,
         \gbuff[15][25] , \gbuff[15][24] , \gbuff[15][23] , \gbuff[15][22] ,
         \gbuff[15][21] , \gbuff[15][20] , \gbuff[15][19] , \gbuff[15][18] ,
         \gbuff[15][17] , \gbuff[15][16] , \gbuff[15][15] , \gbuff[15][14] ,
         \gbuff[15][13] , \gbuff[15][12] , \gbuff[15][11] , \gbuff[15][10] ,
         \gbuff[15][9] , \gbuff[15][8] , \gbuff[15][7] , \gbuff[15][6] ,
         \gbuff[15][5] , \gbuff[15][4] , \gbuff[15][3] , \gbuff[15][2] ,
         \gbuff[15][1] , \gbuff[15][0] , \gbuff[14][31] , \gbuff[14][30] ,
         \gbuff[14][29] , \gbuff[14][28] , \gbuff[14][27] , \gbuff[14][26] ,
         \gbuff[14][25] , \gbuff[14][24] , \gbuff[14][23] , \gbuff[14][22] ,
         \gbuff[14][21] , \gbuff[14][20] , \gbuff[14][19] , \gbuff[14][18] ,
         \gbuff[14][17] , \gbuff[14][16] , \gbuff[14][15] , \gbuff[14][14] ,
         \gbuff[14][13] , \gbuff[14][12] , \gbuff[14][11] , \gbuff[14][10] ,
         \gbuff[14][9] , \gbuff[14][8] , \gbuff[14][7] , \gbuff[14][6] ,
         \gbuff[14][5] , \gbuff[14][4] , \gbuff[14][3] , \gbuff[14][2] ,
         \gbuff[14][1] , \gbuff[14][0] , \gbuff[17][31] , \gbuff[17][30] ,
         \gbuff[17][29] , \gbuff[17][28] , \gbuff[17][27] , \gbuff[17][26] ,
         \gbuff[17][25] , \gbuff[17][24] , \gbuff[17][23] , \gbuff[17][22] ,
         \gbuff[17][21] , \gbuff[17][20] , \gbuff[17][19] , \gbuff[17][18] ,
         \gbuff[17][17] , \gbuff[17][16] , \gbuff[17][15] , \gbuff[17][14] ,
         \gbuff[17][13] , \gbuff[17][12] , \gbuff[17][11] , \gbuff[17][10] ,
         \gbuff[17][9] , \gbuff[17][8] , \gbuff[17][7] , \gbuff[17][6] ,
         \gbuff[17][5] , \gbuff[17][4] , \gbuff[17][3] , \gbuff[17][2] ,
         \gbuff[17][1] , \gbuff[17][0] , \gbuff[16][31] , \gbuff[16][30] ,
         \gbuff[16][29] , \gbuff[16][28] , \gbuff[16][27] , \gbuff[16][26] ,
         \gbuff[16][25] , \gbuff[16][24] , \gbuff[16][23] , \gbuff[16][22] ,
         \gbuff[16][21] , \gbuff[16][20] , \gbuff[16][19] , \gbuff[16][18] ,
         \gbuff[16][17] , \gbuff[16][16] , \gbuff[16][15] , \gbuff[16][14] ,
         \gbuff[16][13] , \gbuff[16][12] , \gbuff[16][11] , \gbuff[16][10] ,
         \gbuff[16][9] , \gbuff[16][8] , \gbuff[16][7] , \gbuff[16][6] ,
         \gbuff[16][5] , \gbuff[16][4] , \gbuff[16][3] , \gbuff[16][2] ,
         \gbuff[16][1] , \gbuff[16][0] , \gbuff[19][31] , \gbuff[19][30] ,
         \gbuff[19][29] , \gbuff[19][28] , \gbuff[19][27] , \gbuff[19][26] ,
         \gbuff[19][25] , \gbuff[19][24] , \gbuff[19][23] , \gbuff[19][22] ,
         \gbuff[19][21] , \gbuff[19][20] , \gbuff[19][19] , \gbuff[19][18] ,
         \gbuff[19][17] , \gbuff[19][16] , \gbuff[19][15] , \gbuff[19][14] ,
         \gbuff[19][13] , \gbuff[19][12] , \gbuff[19][11] , \gbuff[19][10] ,
         \gbuff[19][9] , \gbuff[19][8] , \gbuff[19][7] , \gbuff[19][6] ,
         \gbuff[19][5] , \gbuff[19][4] , \gbuff[19][3] , \gbuff[19][2] ,
         \gbuff[19][1] , \gbuff[19][0] , \gbuff[18][31] , \gbuff[18][30] ,
         \gbuff[18][29] , \gbuff[18][28] , \gbuff[18][27] , \gbuff[18][26] ,
         \gbuff[18][25] , \gbuff[18][24] , \gbuff[18][23] , \gbuff[18][22] ,
         \gbuff[18][21] , \gbuff[18][20] , \gbuff[18][19] , \gbuff[18][18] ,
         \gbuff[18][17] , \gbuff[18][16] , \gbuff[18][15] , \gbuff[18][14] ,
         \gbuff[18][13] , \gbuff[18][12] , \gbuff[18][11] , \gbuff[18][10] ,
         \gbuff[18][9] , \gbuff[18][8] , \gbuff[18][7] , \gbuff[18][6] ,
         \gbuff[18][5] , \gbuff[18][4] , \gbuff[18][3] , \gbuff[18][2] ,
         \gbuff[18][1] , \gbuff[18][0] , \gbuff[21][31] , \gbuff[21][30] ,
         \gbuff[21][29] , \gbuff[21][28] , \gbuff[21][27] , \gbuff[21][26] ,
         \gbuff[21][25] , \gbuff[21][24] , \gbuff[21][23] , \gbuff[21][22] ,
         \gbuff[21][21] , \gbuff[21][20] , \gbuff[21][19] , \gbuff[21][18] ,
         \gbuff[21][17] , \gbuff[21][16] , \gbuff[21][15] , \gbuff[21][14] ,
         \gbuff[21][13] , \gbuff[21][12] , \gbuff[21][11] , \gbuff[21][10] ,
         \gbuff[21][9] , \gbuff[21][8] , \gbuff[21][7] , \gbuff[21][6] ,
         \gbuff[21][5] , \gbuff[21][4] , \gbuff[21][3] , \gbuff[21][2] ,
         \gbuff[21][1] , \gbuff[21][0] , \gbuff[20][31] , \gbuff[20][30] ,
         \gbuff[20][29] , \gbuff[20][28] , \gbuff[20][27] , \gbuff[20][26] ,
         \gbuff[20][25] , \gbuff[20][24] , \gbuff[20][23] , \gbuff[20][22] ,
         \gbuff[20][21] , \gbuff[20][20] , \gbuff[20][19] , \gbuff[20][18] ,
         \gbuff[20][17] , \gbuff[20][16] , \gbuff[20][15] , \gbuff[20][14] ,
         \gbuff[20][13] , \gbuff[20][12] , \gbuff[20][11] , \gbuff[20][10] ,
         \gbuff[20][9] , \gbuff[20][8] , \gbuff[20][7] , \gbuff[20][6] ,
         \gbuff[20][5] , \gbuff[20][4] , \gbuff[20][3] , \gbuff[20][2] ,
         \gbuff[20][1] , \gbuff[20][0] , \gbuff[23][31] , \gbuff[23][30] ,
         \gbuff[23][29] , \gbuff[23][28] , \gbuff[23][27] , \gbuff[23][26] ,
         \gbuff[23][25] , \gbuff[23][24] , \gbuff[23][23] , \gbuff[23][22] ,
         \gbuff[23][21] , \gbuff[23][20] , \gbuff[23][19] , \gbuff[23][18] ,
         \gbuff[23][17] , \gbuff[23][16] , \gbuff[23][15] , \gbuff[23][14] ,
         \gbuff[23][13] , \gbuff[23][12] , \gbuff[23][11] , \gbuff[23][10] ,
         \gbuff[23][9] , \gbuff[23][8] , \gbuff[23][7] , \gbuff[23][6] ,
         \gbuff[23][5] , \gbuff[23][4] , \gbuff[23][3] , \gbuff[23][2] ,
         \gbuff[23][1] , \gbuff[23][0] , \gbuff[22][31] , \gbuff[22][30] ,
         \gbuff[22][29] , \gbuff[22][28] , \gbuff[22][27] , \gbuff[22][26] ,
         \gbuff[22][25] , \gbuff[22][24] , \gbuff[22][23] , \gbuff[22][22] ,
         \gbuff[22][21] , \gbuff[22][20] , \gbuff[22][19] , \gbuff[22][18] ,
         \gbuff[22][17] , \gbuff[22][16] , \gbuff[22][15] , \gbuff[22][14] ,
         \gbuff[22][13] , \gbuff[22][12] , \gbuff[22][11] , \gbuff[22][10] ,
         \gbuff[22][9] , \gbuff[22][8] , \gbuff[22][7] , \gbuff[22][6] ,
         \gbuff[22][5] , \gbuff[22][4] , \gbuff[22][3] , \gbuff[22][2] ,
         \gbuff[22][1] , \gbuff[22][0] , \gbuff[25][31] , \gbuff[25][30] ,
         \gbuff[25][29] , \gbuff[25][28] , \gbuff[25][27] , \gbuff[25][26] ,
         \gbuff[25][25] , \gbuff[25][24] , \gbuff[25][23] , \gbuff[25][22] ,
         \gbuff[25][21] , \gbuff[25][20] , \gbuff[25][19] , \gbuff[25][18] ,
         \gbuff[25][17] , \gbuff[25][16] , \gbuff[25][15] , \gbuff[25][14] ,
         \gbuff[25][13] , \gbuff[25][12] , \gbuff[25][11] , \gbuff[25][10] ,
         \gbuff[25][9] , \gbuff[25][8] , \gbuff[25][7] , \gbuff[25][6] ,
         \gbuff[25][5] , \gbuff[25][4] , \gbuff[25][3] , \gbuff[25][2] ,
         \gbuff[25][1] , \gbuff[25][0] , \gbuff[24][31] , \gbuff[24][30] ,
         \gbuff[24][29] , \gbuff[24][28] , \gbuff[24][27] , \gbuff[24][26] ,
         \gbuff[24][25] , \gbuff[24][24] , \gbuff[24][23] , \gbuff[24][22] ,
         \gbuff[24][21] , \gbuff[24][20] , \gbuff[24][19] , \gbuff[24][18] ,
         \gbuff[24][17] , \gbuff[24][16] , \gbuff[24][15] , \gbuff[24][14] ,
         \gbuff[24][13] , \gbuff[24][12] , \gbuff[24][11] , \gbuff[24][10] ,
         \gbuff[24][9] , \gbuff[24][8] , \gbuff[24][7] , \gbuff[24][6] ,
         \gbuff[24][5] , \gbuff[24][4] , \gbuff[24][3] , \gbuff[24][2] ,
         \gbuff[24][1] , \gbuff[24][0] , \gbuff[27][31] , \gbuff[27][30] ,
         \gbuff[27][29] , \gbuff[27][28] , \gbuff[27][27] , \gbuff[27][26] ,
         \gbuff[27][25] , \gbuff[27][24] , \gbuff[27][23] , \gbuff[27][22] ,
         \gbuff[27][21] , \gbuff[27][20] , \gbuff[27][19] , \gbuff[27][18] ,
         \gbuff[27][17] , \gbuff[27][16] , \gbuff[27][15] , \gbuff[27][14] ,
         \gbuff[27][13] , \gbuff[27][12] , \gbuff[27][11] , \gbuff[27][10] ,
         \gbuff[27][9] , \gbuff[27][8] , \gbuff[27][7] , \gbuff[27][6] ,
         \gbuff[27][5] , \gbuff[27][4] , \gbuff[27][3] , \gbuff[27][2] ,
         \gbuff[27][1] , \gbuff[27][0] , \gbuff[26][31] , \gbuff[26][30] ,
         \gbuff[26][29] , \gbuff[26][28] , \gbuff[26][27] , \gbuff[26][26] ,
         \gbuff[26][25] , \gbuff[26][24] , \gbuff[26][23] , \gbuff[26][22] ,
         \gbuff[26][21] , \gbuff[26][20] , \gbuff[26][19] , \gbuff[26][18] ,
         \gbuff[26][17] , \gbuff[26][16] , \gbuff[26][15] , \gbuff[26][14] ,
         \gbuff[26][13] , \gbuff[26][12] , \gbuff[26][11] , \gbuff[26][10] ,
         \gbuff[26][9] , \gbuff[26][8] , \gbuff[26][7] , \gbuff[26][6] ,
         \gbuff[26][5] , \gbuff[26][4] , \gbuff[26][3] , \gbuff[26][2] ,
         \gbuff[26][1] , \gbuff[26][0] , \gbuff[29][31] , \gbuff[29][30] ,
         \gbuff[29][29] , \gbuff[29][28] , \gbuff[29][27] , \gbuff[29][26] ,
         \gbuff[29][25] , \gbuff[29][24] , \gbuff[29][23] , \gbuff[29][22] ,
         \gbuff[29][21] , \gbuff[29][20] , \gbuff[29][19] , \gbuff[29][18] ,
         \gbuff[29][17] , \gbuff[29][16] , \gbuff[29][15] , \gbuff[29][14] ,
         \gbuff[29][13] , \gbuff[29][12] , \gbuff[29][11] , \gbuff[29][10] ,
         \gbuff[29][9] , \gbuff[29][8] , \gbuff[29][7] , \gbuff[29][6] ,
         \gbuff[29][5] , \gbuff[29][4] , \gbuff[29][3] , \gbuff[29][2] ,
         \gbuff[29][1] , \gbuff[29][0] , \gbuff[28][31] , \gbuff[28][30] ,
         \gbuff[28][29] , \gbuff[28][28] , \gbuff[28][27] , \gbuff[28][26] ,
         \gbuff[28][25] , \gbuff[28][24] , \gbuff[28][23] , \gbuff[28][22] ,
         \gbuff[28][21] , \gbuff[28][20] , \gbuff[28][19] , \gbuff[28][18] ,
         \gbuff[28][17] , \gbuff[28][16] , \gbuff[28][15] , \gbuff[28][14] ,
         \gbuff[28][13] , \gbuff[28][12] , \gbuff[28][11] , \gbuff[28][10] ,
         \gbuff[28][9] , \gbuff[28][8] , \gbuff[28][7] , \gbuff[28][6] ,
         \gbuff[28][5] , \gbuff[28][4] , \gbuff[28][3] , \gbuff[28][2] ,
         \gbuff[28][1] , \gbuff[28][0] , \gbuff[31][31] , \gbuff[31][30] ,
         \gbuff[31][29] , \gbuff[31][28] , \gbuff[31][27] , \gbuff[31][26] ,
         \gbuff[31][25] , \gbuff[31][24] , \gbuff[31][23] , \gbuff[31][22] ,
         \gbuff[31][21] , \gbuff[31][20] , \gbuff[31][19] , \gbuff[31][18] ,
         \gbuff[31][17] , \gbuff[31][16] , \gbuff[31][15] , \gbuff[31][14] ,
         \gbuff[31][13] , \gbuff[31][12] , \gbuff[31][11] , \gbuff[31][10] ,
         \gbuff[31][9] , \gbuff[31][8] , \gbuff[31][7] , \gbuff[31][6] ,
         \gbuff[31][5] , \gbuff[31][4] , \gbuff[31][3] , \gbuff[31][2] ,
         \gbuff[31][1] , \gbuff[31][0] , \gbuff[30][31] , \gbuff[30][30] ,
         \gbuff[30][29] , \gbuff[30][28] , \gbuff[30][27] , \gbuff[30][26] ,
         \gbuff[30][25] , \gbuff[30][24] , \gbuff[30][23] , \gbuff[30][22] ,
         \gbuff[30][21] , \gbuff[30][20] , \gbuff[30][19] , \gbuff[30][18] ,
         \gbuff[30][17] , \gbuff[30][16] , \gbuff[30][15] , \gbuff[30][14] ,
         \gbuff[30][13] , \gbuff[30][12] , \gbuff[30][11] , \gbuff[30][10] ,
         \gbuff[30][9] , \gbuff[30][8] , \gbuff[30][7] , \gbuff[30][6] ,
         \gbuff[30][5] , \gbuff[30][4] , \gbuff[30][3] , \gbuff[30][2] ,
         \gbuff[30][1] , \gbuff[30][0] , N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N81, n102,
         n103, n105, n107, n109, n111, n113, n115, n117, n118, n120, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n104, n106, n108, n110, n112, n114, n116, n119,
         n121, n122, n123, n124, n125, n126, n127, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646;
  assign N10 = index[0];
  assign N11 = index[1];
  assign N12 = index[2];
  assign N13 = index[3];
  assign N14 = index[4];

  DFFRX1 \gbuff_reg[29][31]  ( .D(n1105), .CK(clk), .RN(n23), .Q(
        \gbuff[29][31] ) );
  DFFRX1 \gbuff_reg[29][30]  ( .D(n1104), .CK(clk), .RN(n21), .Q(
        \gbuff[29][30] ) );
  DFFRX1 \gbuff_reg[29][29]  ( .D(n1103), .CK(clk), .RN(n24), .Q(
        \gbuff[29][29] ) );
  DFFRX1 \gbuff_reg[29][28]  ( .D(n1102), .CK(clk), .RN(n20), .Q(
        \gbuff[29][28] ) );
  DFFRX1 \gbuff_reg[29][27]  ( .D(n1101), .CK(clk), .RN(n19), .Q(
        \gbuff[29][27] ) );
  DFFRX1 \gbuff_reg[29][26]  ( .D(n1100), .CK(clk), .RN(n24), .Q(
        \gbuff[29][26] ) );
  DFFRX1 \gbuff_reg[29][25]  ( .D(n1099), .CK(clk), .RN(n20), .Q(
        \gbuff[29][25] ) );
  DFFRX1 \gbuff_reg[29][24]  ( .D(n1098), .CK(clk), .RN(n26), .Q(
        \gbuff[29][24] ) );
  DFFRX1 \gbuff_reg[29][23]  ( .D(n1097), .CK(clk), .RN(n17), .Q(
        \gbuff[29][23] ) );
  DFFRX1 \gbuff_reg[29][22]  ( .D(n1096), .CK(clk), .RN(n25), .Q(
        \gbuff[29][22] ) );
  DFFRX1 \gbuff_reg[29][21]  ( .D(n1095), .CK(clk), .RN(n25), .Q(
        \gbuff[29][21] ) );
  DFFRX1 \gbuff_reg[29][20]  ( .D(n1094), .CK(clk), .RN(n23), .Q(
        \gbuff[29][20] ) );
  DFFRX1 \gbuff_reg[29][19]  ( .D(n1093), .CK(clk), .RN(n19), .Q(
        \gbuff[29][19] ) );
  DFFRX1 \gbuff_reg[29][18]  ( .D(n1092), .CK(clk), .RN(n18), .Q(
        \gbuff[29][18] ) );
  DFFRX1 \gbuff_reg[29][17]  ( .D(n1091), .CK(clk), .RN(n25), .Q(
        \gbuff[29][17] ) );
  DFFRX1 \gbuff_reg[29][16]  ( .D(n1090), .CK(clk), .RN(n26), .Q(
        \gbuff[29][16] ) );
  DFFRX1 \gbuff_reg[29][15]  ( .D(n1089), .CK(clk), .RN(n21), .Q(
        \gbuff[29][15] ) );
  DFFRX1 \gbuff_reg[29][14]  ( .D(n1088), .CK(clk), .RN(n19), .Q(
        \gbuff[29][14] ) );
  DFFRX1 \gbuff_reg[29][13]  ( .D(n1087), .CK(clk), .RN(n25), .Q(
        \gbuff[29][13] ) );
  DFFRX1 \gbuff_reg[29][12]  ( .D(n1086), .CK(clk), .RN(n23), .Q(
        \gbuff[29][12] ) );
  DFFRX1 \gbuff_reg[29][11]  ( .D(n1085), .CK(clk), .RN(n24), .Q(
        \gbuff[29][11] ) );
  DFFRX1 \gbuff_reg[29][10]  ( .D(n1084), .CK(clk), .RN(n23), .Q(
        \gbuff[29][10] ) );
  DFFRX1 \gbuff_reg[29][9]  ( .D(n1083), .CK(clk), .RN(n21), .Q(\gbuff[29][9] ) );
  DFFRX1 \gbuff_reg[29][8]  ( .D(n1082), .CK(clk), .RN(n20), .Q(\gbuff[29][8] ) );
  DFFRX1 \gbuff_reg[29][7]  ( .D(n1081), .CK(clk), .RN(n21), .Q(\gbuff[29][7] ) );
  DFFRX1 \gbuff_reg[29][6]  ( .D(n1080), .CK(clk), .RN(n19), .Q(\gbuff[29][6] ) );
  DFFRX1 \gbuff_reg[29][5]  ( .D(n1079), .CK(clk), .RN(n17), .Q(\gbuff[29][5] ) );
  DFFRX1 \gbuff_reg[29][4]  ( .D(n1078), .CK(clk), .RN(n18), .Q(\gbuff[29][4] ) );
  DFFRX1 \gbuff_reg[29][3]  ( .D(n1077), .CK(clk), .RN(n20), .Q(\gbuff[29][3] ) );
  DFFRX1 \gbuff_reg[29][2]  ( .D(n1076), .CK(clk), .RN(n25), .Q(\gbuff[29][2] ) );
  DFFRX1 \gbuff_reg[29][1]  ( .D(n1075), .CK(clk), .RN(n24), .Q(\gbuff[29][1] ) );
  DFFRX1 \gbuff_reg[29][0]  ( .D(n1074), .CK(clk), .RN(n24), .Q(\gbuff[29][0] ) );
  DFFRX1 \gbuff_reg[25][31]  ( .D(n977), .CK(clk), .RN(n26), .Q(
        \gbuff[25][31] ) );
  DFFRX1 \gbuff_reg[25][30]  ( .D(n976), .CK(clk), .RN(n26), .Q(
        \gbuff[25][30] ) );
  DFFRX1 \gbuff_reg[25][29]  ( .D(n975), .CK(clk), .RN(n26), .Q(
        \gbuff[25][29] ) );
  DFFRX1 \gbuff_reg[25][28]  ( .D(n974), .CK(clk), .RN(n19), .Q(
        \gbuff[25][28] ) );
  DFFRX1 \gbuff_reg[25][27]  ( .D(n973), .CK(clk), .RN(n20), .Q(
        \gbuff[25][27] ) );
  DFFRX1 \gbuff_reg[25][26]  ( .D(n972), .CK(clk), .RN(n17), .Q(
        \gbuff[25][26] ) );
  DFFRX1 \gbuff_reg[25][25]  ( .D(n971), .CK(clk), .RN(n23), .Q(
        \gbuff[25][25] ) );
  DFFRX1 \gbuff_reg[25][24]  ( .D(n970), .CK(clk), .RN(n24), .Q(
        \gbuff[25][24] ) );
  DFFRX1 \gbuff_reg[25][23]  ( .D(n969), .CK(clk), .RN(n18), .Q(
        \gbuff[25][23] ) );
  DFFRX1 \gbuff_reg[25][22]  ( .D(n968), .CK(clk), .RN(n23), .Q(
        \gbuff[25][22] ) );
  DFFRX1 \gbuff_reg[25][21]  ( .D(n967), .CK(clk), .RN(n26), .Q(
        \gbuff[25][21] ) );
  DFFRX1 \gbuff_reg[25][20]  ( .D(n966), .CK(clk), .RN(n19), .Q(
        \gbuff[25][20] ) );
  DFFRX1 \gbuff_reg[25][19]  ( .D(n965), .CK(clk), .RN(n25), .Q(
        \gbuff[25][19] ) );
  DFFRX1 \gbuff_reg[25][18]  ( .D(n964), .CK(clk), .RN(n24), .Q(
        \gbuff[25][18] ) );
  DFFRX1 \gbuff_reg[25][17]  ( .D(n963), .CK(clk), .RN(n23), .Q(
        \gbuff[25][17] ) );
  DFFRX1 \gbuff_reg[25][16]  ( .D(n962), .CK(clk), .RN(n21), .Q(
        \gbuff[25][16] ) );
  DFFRX1 \gbuff_reg[25][15]  ( .D(n961), .CK(clk), .RN(n18), .Q(
        \gbuff[25][15] ) );
  DFFRX1 \gbuff_reg[25][14]  ( .D(n960), .CK(clk), .RN(n23), .Q(
        \gbuff[25][14] ) );
  DFFRX1 \gbuff_reg[25][13]  ( .D(n959), .CK(clk), .RN(n18), .Q(
        \gbuff[25][13] ) );
  DFFRX1 \gbuff_reg[25][12]  ( .D(n958), .CK(clk), .RN(n21), .Q(
        \gbuff[25][12] ) );
  DFFRX1 \gbuff_reg[25][11]  ( .D(n957), .CK(clk), .RN(n17), .Q(
        \gbuff[25][11] ) );
  DFFRX1 \gbuff_reg[25][10]  ( .D(n956), .CK(clk), .RN(n17), .Q(
        \gbuff[25][10] ) );
  DFFRX1 \gbuff_reg[25][9]  ( .D(n955), .CK(clk), .RN(n21), .Q(\gbuff[25][9] )
         );
  DFFRX1 \gbuff_reg[25][8]  ( .D(n954), .CK(clk), .RN(n17), .Q(\gbuff[25][8] )
         );
  DFFRX1 \gbuff_reg[25][7]  ( .D(n953), .CK(clk), .RN(n23), .Q(\gbuff[25][7] )
         );
  DFFRX1 \gbuff_reg[25][6]  ( .D(n952), .CK(clk), .RN(n24), .Q(\gbuff[25][6] )
         );
  DFFRX1 \gbuff_reg[25][5]  ( .D(n951), .CK(clk), .RN(n24), .Q(\gbuff[25][5] )
         );
  DFFRX1 \gbuff_reg[25][4]  ( .D(n950), .CK(clk), .RN(n21), .Q(\gbuff[25][4] )
         );
  DFFRX1 \gbuff_reg[25][3]  ( .D(n949), .CK(clk), .RN(n17), .Q(\gbuff[25][3] )
         );
  DFFRX1 \gbuff_reg[25][2]  ( .D(n948), .CK(clk), .RN(n24), .Q(\gbuff[25][2] )
         );
  DFFRX1 \gbuff_reg[25][1]  ( .D(n947), .CK(clk), .RN(n19), .Q(\gbuff[25][1] )
         );
  DFFRX1 \gbuff_reg[25][0]  ( .D(n946), .CK(clk), .RN(n17), .Q(\gbuff[25][0] )
         );
  DFFRX1 \gbuff_reg[21][31]  ( .D(n849), .CK(clk), .RN(n24), .Q(
        \gbuff[21][31] ) );
  DFFRX1 \gbuff_reg[21][30]  ( .D(n848), .CK(clk), .RN(n25), .Q(
        \gbuff[21][30] ) );
  DFFRX1 \gbuff_reg[21][29]  ( .D(n847), .CK(clk), .RN(n24), .Q(
        \gbuff[21][29] ) );
  DFFRX1 \gbuff_reg[21][28]  ( .D(n846), .CK(clk), .RN(n25), .Q(
        \gbuff[21][28] ) );
  DFFRX1 \gbuff_reg[21][27]  ( .D(n845), .CK(clk), .RN(n19), .Q(
        \gbuff[21][27] ) );
  DFFRX1 \gbuff_reg[21][26]  ( .D(n844), .CK(clk), .RN(n25), .Q(
        \gbuff[21][26] ) );
  DFFRX1 \gbuff_reg[21][25]  ( .D(n843), .CK(clk), .RN(n19), .Q(
        \gbuff[21][25] ) );
  DFFRX1 \gbuff_reg[21][24]  ( .D(n842), .CK(clk), .RN(n19), .Q(
        \gbuff[21][24] ) );
  DFFRX1 \gbuff_reg[21][23]  ( .D(n841), .CK(clk), .RN(n24), .Q(
        \gbuff[21][23] ) );
  DFFRX1 \gbuff_reg[21][22]  ( .D(n840), .CK(clk), .RN(n25), .Q(
        \gbuff[21][22] ) );
  DFFRX1 \gbuff_reg[21][21]  ( .D(n839), .CK(clk), .RN(n20), .Q(
        \gbuff[21][21] ) );
  DFFRX1 \gbuff_reg[21][20]  ( .D(n838), .CK(clk), .RN(n20), .Q(
        \gbuff[21][20] ) );
  DFFRX1 \gbuff_reg[21][19]  ( .D(n837), .CK(clk), .RN(n26), .Q(
        \gbuff[21][19] ) );
  DFFRX1 \gbuff_reg[21][18]  ( .D(n836), .CK(clk), .RN(n26), .Q(
        \gbuff[21][18] ) );
  DFFRX1 \gbuff_reg[21][17]  ( .D(n835), .CK(clk), .RN(n17), .Q(
        \gbuff[21][17] ) );
  DFFRX1 \gbuff_reg[21][16]  ( .D(n834), .CK(clk), .RN(n18), .Q(
        \gbuff[21][16] ) );
  DFFRX1 \gbuff_reg[21][15]  ( .D(n833), .CK(clk), .RN(n21), .Q(
        \gbuff[21][15] ) );
  DFFRX1 \gbuff_reg[21][14]  ( .D(n832), .CK(clk), .RN(n17), .Q(
        \gbuff[21][14] ) );
  DFFRX1 \gbuff_reg[21][13]  ( .D(n831), .CK(clk), .RN(n17), .Q(
        \gbuff[21][13] ) );
  DFFRX1 \gbuff_reg[21][12]  ( .D(n830), .CK(clk), .RN(n20), .Q(
        \gbuff[21][12] ) );
  DFFRX1 \gbuff_reg[21][11]  ( .D(n829), .CK(clk), .RN(n26), .Q(
        \gbuff[21][11] ) );
  DFFRX1 \gbuff_reg[21][10]  ( .D(n828), .CK(clk), .RN(n26), .Q(
        \gbuff[21][10] ) );
  DFFRX1 \gbuff_reg[21][9]  ( .D(n827), .CK(clk), .RN(n21), .Q(\gbuff[21][9] )
         );
  DFFRX1 \gbuff_reg[21][8]  ( .D(n826), .CK(clk), .RN(n18), .Q(\gbuff[21][8] )
         );
  DFFRX1 \gbuff_reg[21][7]  ( .D(n825), .CK(clk), .RN(n25), .Q(\gbuff[21][7] )
         );
  DFFRX1 \gbuff_reg[21][6]  ( .D(n824), .CK(clk), .RN(n26), .Q(\gbuff[21][6] )
         );
  DFFRX1 \gbuff_reg[21][5]  ( .D(n823), .CK(clk), .RN(n17), .Q(\gbuff[21][5] )
         );
  DFFRX1 \gbuff_reg[21][4]  ( .D(n822), .CK(clk), .RN(n23), .Q(\gbuff[21][4] )
         );
  DFFRX1 \gbuff_reg[21][3]  ( .D(n821), .CK(clk), .RN(n20), .Q(\gbuff[21][3] )
         );
  DFFRX1 \gbuff_reg[21][2]  ( .D(n820), .CK(clk), .RN(n17), .Q(\gbuff[21][2] )
         );
  DFFRX1 \gbuff_reg[21][1]  ( .D(n819), .CK(clk), .RN(n25), .Q(\gbuff[21][1] )
         );
  DFFRX1 \gbuff_reg[21][0]  ( .D(n818), .CK(clk), .RN(n23), .Q(\gbuff[21][0] )
         );
  DFFRX1 \gbuff_reg[17][31]  ( .D(n721), .CK(clk), .RN(n25), .Q(
        \gbuff[17][31] ) );
  DFFRX1 \gbuff_reg[17][30]  ( .D(n720), .CK(clk), .RN(n26), .Q(
        \gbuff[17][30] ) );
  DFFRX1 \gbuff_reg[17][29]  ( .D(n719), .CK(clk), .RN(n21), .Q(
        \gbuff[17][29] ) );
  DFFRX1 \gbuff_reg[17][28]  ( .D(n718), .CK(clk), .RN(n19), .Q(
        \gbuff[17][28] ) );
  DFFRX1 \gbuff_reg[17][27]  ( .D(n717), .CK(clk), .RN(n23), .Q(
        \gbuff[17][27] ) );
  DFFRX1 \gbuff_reg[17][26]  ( .D(n716), .CK(clk), .RN(n18), .Q(
        \gbuff[17][26] ) );
  DFFRX1 \gbuff_reg[17][25]  ( .D(n715), .CK(clk), .RN(n19), .Q(
        \gbuff[17][25] ) );
  DFFRX1 \gbuff_reg[17][24]  ( .D(n714), .CK(clk), .RN(n20), .Q(
        \gbuff[17][24] ) );
  DFFRX1 \gbuff_reg[17][23]  ( .D(n713), .CK(clk), .RN(n18), .Q(
        \gbuff[17][23] ) );
  DFFRX1 \gbuff_reg[17][22]  ( .D(n712), .CK(clk), .RN(n18), .Q(
        \gbuff[17][22] ) );
  DFFRX1 \gbuff_reg[17][21]  ( .D(n711), .CK(clk), .RN(n18), .Q(
        \gbuff[17][21] ) );
  DFFRX1 \gbuff_reg[17][20]  ( .D(n710), .CK(clk), .RN(n18), .Q(
        \gbuff[17][20] ) );
  DFFRX1 \gbuff_reg[17][19]  ( .D(n709), .CK(clk), .RN(n23), .Q(
        \gbuff[17][19] ) );
  DFFRX1 \gbuff_reg[17][18]  ( .D(n708), .CK(clk), .RN(n25), .Q(
        \gbuff[17][18] ) );
  DFFRX1 \gbuff_reg[17][17]  ( .D(n707), .CK(clk), .RN(n20), .Q(
        \gbuff[17][17] ) );
  DFFRX1 \gbuff_reg[17][16]  ( .D(n706), .CK(clk), .RN(n20), .Q(
        \gbuff[17][16] ) );
  DFFRX1 \gbuff_reg[17][15]  ( .D(n705), .CK(clk), .RN(n19), .Q(
        \gbuff[17][15] ) );
  DFFRX1 \gbuff_reg[17][14]  ( .D(n704), .CK(clk), .RN(n24), .Q(
        \gbuff[17][14] ) );
  DFFRX1 \gbuff_reg[17][13]  ( .D(n703), .CK(clk), .RN(n18), .Q(
        \gbuff[17][13] ) );
  DFFRX1 \gbuff_reg[17][12]  ( .D(n702), .CK(clk), .RN(n26), .Q(
        \gbuff[17][12] ) );
  DFFRX1 \gbuff_reg[17][11]  ( .D(n701), .CK(clk), .RN(n17), .Q(
        \gbuff[17][11] ) );
  DFFRX1 \gbuff_reg[17][10]  ( .D(n700), .CK(clk), .RN(n26), .Q(
        \gbuff[17][10] ) );
  DFFRX1 \gbuff_reg[17][9]  ( .D(n699), .CK(clk), .RN(n23), .Q(\gbuff[17][9] )
         );
  DFFRX1 \gbuff_reg[17][8]  ( .D(n698), .CK(clk), .RN(n25), .Q(\gbuff[17][8] )
         );
  DFFRX1 \gbuff_reg[17][7]  ( .D(n697), .CK(clk), .RN(n19), .Q(\gbuff[17][7] )
         );
  DFFRX1 \gbuff_reg[17][6]  ( .D(n696), .CK(clk), .RN(n24), .Q(\gbuff[17][6] )
         );
  DFFRX1 \gbuff_reg[17][5]  ( .D(n695), .CK(clk), .RN(n19), .Q(\gbuff[17][5] )
         );
  DFFRX1 \gbuff_reg[17][4]  ( .D(n694), .CK(clk), .RN(n21), .Q(\gbuff[17][4] )
         );
  DFFRX1 \gbuff_reg[17][3]  ( .D(n693), .CK(clk), .RN(n21), .Q(\gbuff[17][3] )
         );
  DFFRX1 \gbuff_reg[17][2]  ( .D(n692), .CK(clk), .RN(n24), .Q(\gbuff[17][2] )
         );
  DFFRX1 \gbuff_reg[17][1]  ( .D(n691), .CK(clk), .RN(n18), .Q(\gbuff[17][1] )
         );
  DFFRX1 \gbuff_reg[17][0]  ( .D(n690), .CK(clk), .RN(n21), .Q(\gbuff[17][0] )
         );
  DFFRX1 \gbuff_reg[13][31]  ( .D(n593), .CK(clk), .RN(n24), .Q(
        \gbuff[13][31] ) );
  DFFRX1 \gbuff_reg[13][30]  ( .D(n592), .CK(clk), .RN(n20), .Q(
        \gbuff[13][30] ) );
  DFFRX1 \gbuff_reg[13][29]  ( .D(n591), .CK(clk), .RN(n20), .Q(
        \gbuff[13][29] ) );
  DFFRX1 \gbuff_reg[13][28]  ( .D(n590), .CK(clk), .RN(n17), .Q(
        \gbuff[13][28] ) );
  DFFRX1 \gbuff_reg[13][27]  ( .D(n589), .CK(clk), .RN(n21), .Q(
        \gbuff[13][27] ) );
  DFFRX1 \gbuff_reg[13][26]  ( .D(n588), .CK(clk), .RN(n23), .Q(
        \gbuff[13][26] ) );
  DFFRX1 \gbuff_reg[13][25]  ( .D(n587), .CK(clk), .RN(n18), .Q(
        \gbuff[13][25] ) );
  DFFRX1 \gbuff_reg[13][24]  ( .D(n586), .CK(clk), .RN(n21), .Q(
        \gbuff[13][24] ) );
  DFFRX1 \gbuff_reg[13][23]  ( .D(n585), .CK(clk), .RN(n20), .Q(
        \gbuff[13][23] ) );
  DFFRX1 \gbuff_reg[13][22]  ( .D(n584), .CK(clk), .RN(n17), .Q(
        \gbuff[13][22] ) );
  DFFRX1 \gbuff_reg[13][21]  ( .D(n583), .CK(clk), .RN(n20), .Q(
        \gbuff[13][21] ) );
  DFFRX1 \gbuff_reg[13][20]  ( .D(n582), .CK(clk), .RN(n25), .Q(
        \gbuff[13][20] ) );
  DFFRX1 \gbuff_reg[13][19]  ( .D(n581), .CK(clk), .RN(n26), .Q(
        \gbuff[13][19] ) );
  DFFRX1 \gbuff_reg[13][18]  ( .D(n580), .CK(clk), .RN(n18), .Q(
        \gbuff[13][18] ) );
  DFFRX1 \gbuff_reg[13][17]  ( .D(n579), .CK(clk), .RN(n26), .Q(
        \gbuff[13][17] ) );
  DFFRX1 \gbuff_reg[13][16]  ( .D(n578), .CK(clk), .RN(n26), .Q(
        \gbuff[13][16] ) );
  DFFRX1 \gbuff_reg[13][15]  ( .D(n577), .CK(clk), .RN(n20), .Q(
        \gbuff[13][15] ) );
  DFFRX1 \gbuff_reg[13][14]  ( .D(n576), .CK(clk), .RN(n17), .Q(
        \gbuff[13][14] ) );
  DFFRX1 \gbuff_reg[13][13]  ( .D(n575), .CK(clk), .RN(n23), .Q(
        \gbuff[13][13] ) );
  DFFRX1 \gbuff_reg[13][12]  ( .D(n574), .CK(clk), .RN(n23), .Q(
        \gbuff[13][12] ) );
  DFFRX1 \gbuff_reg[13][11]  ( .D(n573), .CK(clk), .RN(n18), .Q(
        \gbuff[13][11] ) );
  DFFRX1 \gbuff_reg[13][10]  ( .D(n572), .CK(clk), .RN(n20), .Q(
        \gbuff[13][10] ) );
  DFFRX1 \gbuff_reg[13][9]  ( .D(n571), .CK(clk), .RN(n23), .Q(\gbuff[13][9] )
         );
  DFFRX1 \gbuff_reg[13][8]  ( .D(n570), .CK(clk), .RN(n19), .Q(\gbuff[13][8] )
         );
  DFFRX1 \gbuff_reg[13][7]  ( .D(n569), .CK(clk), .RN(n25), .Q(\gbuff[13][7] )
         );
  DFFRX1 \gbuff_reg[13][6]  ( .D(n568), .CK(clk), .RN(n21), .Q(\gbuff[13][6] )
         );
  DFFRX1 \gbuff_reg[13][5]  ( .D(n567), .CK(clk), .RN(n21), .Q(\gbuff[13][5] )
         );
  DFFRX1 \gbuff_reg[13][4]  ( .D(n566), .CK(clk), .RN(n24), .Q(\gbuff[13][4] )
         );
  DFFRX1 \gbuff_reg[13][3]  ( .D(n565), .CK(clk), .RN(n18), .Q(\gbuff[13][3] )
         );
  DFFRX1 \gbuff_reg[13][2]  ( .D(n564), .CK(clk), .RN(n19), .Q(\gbuff[13][2] )
         );
  DFFRX1 \gbuff_reg[13][1]  ( .D(n563), .CK(clk), .RN(n17), .Q(\gbuff[13][1] )
         );
  DFFRX1 \gbuff_reg[13][0]  ( .D(n562), .CK(clk), .RN(n19), .Q(\gbuff[13][0] )
         );
  DFFRX1 \gbuff_reg[9][31]  ( .D(n465), .CK(clk), .RN(n17), .Q(\gbuff[9][31] )
         );
  DFFRX1 \gbuff_reg[9][30]  ( .D(n464), .CK(clk), .RN(n18), .Q(\gbuff[9][30] )
         );
  DFFRX1 \gbuff_reg[9][29]  ( .D(n463), .CK(clk), .RN(n21), .Q(\gbuff[9][29] )
         );
  DFFRX1 \gbuff_reg[9][28]  ( .D(n462), .CK(clk), .RN(n24), .Q(\gbuff[9][28] )
         );
  DFFRX1 \gbuff_reg[9][27]  ( .D(n461), .CK(clk), .RN(n23), .Q(\gbuff[9][27] )
         );
  DFFRX1 \gbuff_reg[9][26]  ( .D(n460), .CK(clk), .RN(n24), .Q(\gbuff[9][26] )
         );
  DFFRX1 \gbuff_reg[9][25]  ( .D(n459), .CK(clk), .RN(n25), .Q(\gbuff[9][25] )
         );
  DFFRX1 \gbuff_reg[9][24]  ( .D(n458), .CK(clk), .RN(n24), .Q(\gbuff[9][24] )
         );
  DFFRX1 \gbuff_reg[9][23]  ( .D(n457), .CK(clk), .RN(n17), .Q(\gbuff[9][23] )
         );
  DFFRX1 \gbuff_reg[9][22]  ( .D(n456), .CK(clk), .RN(n18), .Q(\gbuff[9][22] )
         );
  DFFRX1 \gbuff_reg[9][21]  ( .D(n455), .CK(clk), .RN(n25), .Q(\gbuff[9][21] )
         );
  DFFRX1 \gbuff_reg[9][20]  ( .D(n454), .CK(clk), .RN(n19), .Q(\gbuff[9][20] )
         );
  DFFRX1 \gbuff_reg[9][19]  ( .D(n453), .CK(clk), .RN(n24), .Q(\gbuff[9][19] )
         );
  DFFRX1 \gbuff_reg[9][18]  ( .D(n452), .CK(clk), .RN(n17), .Q(\gbuff[9][18] )
         );
  DFFRX1 \gbuff_reg[9][17]  ( .D(n451), .CK(clk), .RN(n20), .Q(\gbuff[9][17] )
         );
  DFFRX1 \gbuff_reg[9][16]  ( .D(n450), .CK(clk), .RN(n23), .Q(\gbuff[9][16] )
         );
  DFFRX1 \gbuff_reg[9][15]  ( .D(n449), .CK(clk), .RN(n19), .Q(\gbuff[9][15] )
         );
  DFFRX1 \gbuff_reg[9][14]  ( .D(n448), .CK(clk), .RN(n19), .Q(\gbuff[9][14] )
         );
  DFFRX1 \gbuff_reg[9][13]  ( .D(n447), .CK(clk), .RN(n19), .Q(\gbuff[9][13] )
         );
  DFFRX1 \gbuff_reg[9][12]  ( .D(n446), .CK(clk), .RN(n26), .Q(\gbuff[9][12] )
         );
  DFFRX1 \gbuff_reg[9][11]  ( .D(n445), .CK(clk), .RN(n24), .Q(\gbuff[9][11] )
         );
  DFFRX1 \gbuff_reg[9][10]  ( .D(n444), .CK(clk), .RN(n21), .Q(\gbuff[9][10] )
         );
  DFFRX1 \gbuff_reg[9][9]  ( .D(n443), .CK(clk), .RN(n24), .Q(\gbuff[9][9] )
         );
  DFFRX1 \gbuff_reg[9][8]  ( .D(n442), .CK(clk), .RN(n23), .Q(\gbuff[9][8] )
         );
  DFFRX1 \gbuff_reg[9][7]  ( .D(n441), .CK(clk), .RN(n26), .Q(\gbuff[9][7] )
         );
  DFFRX1 \gbuff_reg[9][6]  ( .D(n440), .CK(clk), .RN(n20), .Q(\gbuff[9][6] )
         );
  DFFRX1 \gbuff_reg[9][5]  ( .D(n439), .CK(clk), .RN(n19), .Q(\gbuff[9][5] )
         );
  DFFRX1 \gbuff_reg[9][4]  ( .D(n438), .CK(clk), .RN(n26), .Q(\gbuff[9][4] )
         );
  DFFRX1 \gbuff_reg[9][3]  ( .D(n437), .CK(clk), .RN(n21), .Q(\gbuff[9][3] )
         );
  DFFRX1 \gbuff_reg[9][2]  ( .D(n436), .CK(clk), .RN(n20), .Q(\gbuff[9][2] )
         );
  DFFRX1 \gbuff_reg[9][1]  ( .D(n435), .CK(clk), .RN(n24), .Q(\gbuff[9][1] )
         );
  DFFRX1 \gbuff_reg[9][0]  ( .D(n434), .CK(clk), .RN(n17), .Q(\gbuff[9][0] )
         );
  DFFRX1 \gbuff_reg[5][31]  ( .D(n337), .CK(clk), .RN(n26), .Q(\gbuff[5][31] )
         );
  DFFRX1 \gbuff_reg[5][30]  ( .D(n336), .CK(clk), .RN(n20), .Q(\gbuff[5][30] )
         );
  DFFRX1 \gbuff_reg[5][29]  ( .D(n335), .CK(clk), .RN(n26), .Q(\gbuff[5][29] )
         );
  DFFRX1 \gbuff_reg[5][28]  ( .D(n334), .CK(clk), .RN(n25), .Q(\gbuff[5][28] )
         );
  DFFRX1 \gbuff_reg[5][27]  ( .D(n333), .CK(clk), .RN(n25), .Q(\gbuff[5][27] )
         );
  DFFRX1 \gbuff_reg[5][26]  ( .D(n332), .CK(clk), .RN(n21), .Q(\gbuff[5][26] )
         );
  DFFRX1 \gbuff_reg[5][25]  ( .D(n331), .CK(clk), .RN(n25), .Q(\gbuff[5][25] )
         );
  DFFRX1 \gbuff_reg[5][24]  ( .D(n330), .CK(clk), .RN(n25), .Q(\gbuff[5][24] )
         );
  DFFRX1 \gbuff_reg[5][23]  ( .D(n329), .CK(clk), .RN(n20), .Q(\gbuff[5][23] )
         );
  DFFRX1 \gbuff_reg[5][22]  ( .D(n328), .CK(clk), .RN(n23), .Q(\gbuff[5][22] )
         );
  DFFRX1 \gbuff_reg[5][21]  ( .D(n327), .CK(clk), .RN(n23), .Q(\gbuff[5][21] )
         );
  DFFRX1 \gbuff_reg[5][20]  ( .D(n326), .CK(clk), .RN(n25), .Q(\gbuff[5][20] )
         );
  DFFRX1 \gbuff_reg[5][19]  ( .D(n325), .CK(clk), .RN(n25), .Q(\gbuff[5][19] )
         );
  DFFRX1 \gbuff_reg[5][18]  ( .D(n324), .CK(clk), .RN(n20), .Q(\gbuff[5][18] )
         );
  DFFRX1 \gbuff_reg[5][17]  ( .D(n323), .CK(clk), .RN(n26), .Q(\gbuff[5][17] )
         );
  DFFRX1 \gbuff_reg[5][16]  ( .D(n322), .CK(clk), .RN(n25), .Q(\gbuff[5][16] )
         );
  DFFRX1 \gbuff_reg[5][15]  ( .D(n321), .CK(clk), .RN(n23), .Q(\gbuff[5][15] )
         );
  DFFRX1 \gbuff_reg[5][14]  ( .D(n320), .CK(clk), .RN(n21), .Q(\gbuff[5][14] )
         );
  DFFRX1 \gbuff_reg[5][13]  ( .D(n319), .CK(clk), .RN(n23), .Q(\gbuff[5][13] )
         );
  DFFRX1 \gbuff_reg[5][12]  ( .D(n318), .CK(clk), .RN(n17), .Q(\gbuff[5][12] )
         );
  DFFRX1 \gbuff_reg[5][11]  ( .D(n317), .CK(clk), .RN(n18), .Q(\gbuff[5][11] )
         );
  DFFRX1 \gbuff_reg[5][10]  ( .D(n316), .CK(clk), .RN(n17), .Q(\gbuff[5][10] )
         );
  DFFRX1 \gbuff_reg[5][9]  ( .D(n315), .CK(clk), .RN(n26), .Q(\gbuff[5][9] )
         );
  DFFRX1 \gbuff_reg[5][8]  ( .D(n314), .CK(clk), .RN(n18), .Q(\gbuff[5][8] )
         );
  DFFRX1 \gbuff_reg[5][7]  ( .D(n313), .CK(clk), .RN(n23), .Q(\gbuff[5][7] )
         );
  DFFRX1 \gbuff_reg[5][6]  ( .D(n312), .CK(clk), .RN(n21), .Q(\gbuff[5][6] )
         );
  DFFRX1 \gbuff_reg[5][5]  ( .D(n311), .CK(clk), .RN(n24), .Q(\gbuff[5][5] )
         );
  DFFRX1 \gbuff_reg[5][4]  ( .D(n310), .CK(clk), .RN(n23), .Q(\gbuff[5][4] )
         );
  DFFRX1 \gbuff_reg[5][3]  ( .D(n309), .CK(clk), .RN(n19), .Q(\gbuff[5][3] )
         );
  DFFRX1 \gbuff_reg[5][2]  ( .D(n308), .CK(clk), .RN(n18), .Q(\gbuff[5][2] )
         );
  DFFRX1 \gbuff_reg[5][1]  ( .D(n307), .CK(clk), .RN(n21), .Q(\gbuff[5][1] )
         );
  DFFRX1 \gbuff_reg[5][0]  ( .D(n306), .CK(clk), .RN(n26), .Q(\gbuff[5][0] )
         );
  DFFRX1 \gbuff_reg[1][31]  ( .D(n209), .CK(clk), .RN(n17), .Q(\gbuff[1][31] )
         );
  DFFRX1 \gbuff_reg[1][30]  ( .D(n208), .CK(clk), .RN(n25), .Q(\gbuff[1][30] )
         );
  DFFRX1 \gbuff_reg[1][29]  ( .D(n207), .CK(clk), .RN(n25), .Q(\gbuff[1][29] )
         );
  DFFRX1 \gbuff_reg[1][28]  ( .D(n206), .CK(clk), .RN(n23), .Q(\gbuff[1][28] )
         );
  DFFRX1 \gbuff_reg[1][27]  ( .D(n205), .CK(clk), .RN(n19), .Q(\gbuff[1][27] )
         );
  DFFRX1 \gbuff_reg[1][26]  ( .D(n204), .CK(clk), .RN(n18), .Q(\gbuff[1][26] )
         );
  DFFRX1 \gbuff_reg[1][25]  ( .D(n203), .CK(clk), .RN(n25), .Q(\gbuff[1][25] )
         );
  DFFRX1 \gbuff_reg[1][24]  ( .D(n202), .CK(clk), .RN(n26), .Q(\gbuff[1][24] )
         );
  DFFRX1 \gbuff_reg[1][23]  ( .D(n201), .CK(clk), .RN(n21), .Q(\gbuff[1][23] )
         );
  DFFRX1 \gbuff_reg[1][22]  ( .D(n200), .CK(clk), .RN(n19), .Q(\gbuff[1][22] )
         );
  DFFRX1 \gbuff_reg[1][21]  ( .D(n199), .CK(clk), .RN(n25), .Q(\gbuff[1][21] )
         );
  DFFRX1 \gbuff_reg[1][20]  ( .D(n198), .CK(clk), .RN(n24), .Q(\gbuff[1][20] )
         );
  DFFRX1 \gbuff_reg[1][19]  ( .D(n197), .CK(clk), .RN(n24), .Q(\gbuff[1][19] )
         );
  DFFRX1 \gbuff_reg[1][18]  ( .D(n196), .CK(clk), .RN(n21), .Q(\gbuff[1][18] )
         );
  DFFRX1 \gbuff_reg[1][17]  ( .D(n195), .CK(clk), .RN(n17), .Q(\gbuff[1][17] )
         );
  DFFRX1 \gbuff_reg[1][16]  ( .D(n194), .CK(clk), .RN(n20), .Q(\gbuff[1][16] )
         );
  DFFRX1 \gbuff_reg[1][15]  ( .D(n193), .CK(clk), .RN(n21), .Q(\gbuff[1][15] )
         );
  DFFRX1 \gbuff_reg[1][14]  ( .D(n192), .CK(clk), .RN(n19), .Q(\gbuff[1][14] )
         );
  DFFRX1 \gbuff_reg[1][13]  ( .D(n191), .CK(clk), .RN(n17), .Q(\gbuff[1][13] )
         );
  DFFRX1 \gbuff_reg[1][12]  ( .D(n190), .CK(clk), .RN(n26), .Q(\gbuff[1][12] )
         );
  DFFRX1 \gbuff_reg[1][11]  ( .D(n189), .CK(clk), .RN(n20), .Q(\gbuff[1][11] )
         );
  DFFRX1 \gbuff_reg[1][10]  ( .D(n188), .CK(clk), .RN(n19), .Q(\gbuff[1][10] )
         );
  DFFRX1 \gbuff_reg[1][9]  ( .D(n187), .CK(clk), .RN(n26), .Q(\gbuff[1][9] )
         );
  DFFRX1 \gbuff_reg[1][8]  ( .D(n186), .CK(clk), .RN(n24), .Q(\gbuff[1][8] )
         );
  DFFRX1 \gbuff_reg[1][7]  ( .D(n185), .CK(clk), .RN(n26), .Q(\gbuff[1][7] )
         );
  DFFRX1 \gbuff_reg[1][6]  ( .D(n184), .CK(clk), .RN(n26), .Q(\gbuff[1][6] )
         );
  DFFRX1 \gbuff_reg[1][5]  ( .D(n183), .CK(clk), .RN(n26), .Q(\gbuff[1][5] )
         );
  DFFRX1 \gbuff_reg[1][4]  ( .D(n182), .CK(clk), .RN(n19), .Q(\gbuff[1][4] )
         );
  DFFRX1 \gbuff_reg[1][3]  ( .D(n181), .CK(clk), .RN(n20), .Q(\gbuff[1][3] )
         );
  DFFRX1 \gbuff_reg[1][2]  ( .D(n180), .CK(clk), .RN(n17), .Q(\gbuff[1][2] )
         );
  DFFRX1 \gbuff_reg[1][1]  ( .D(n179), .CK(clk), .RN(n23), .Q(\gbuff[1][1] )
         );
  DFFRX1 \gbuff_reg[1][0]  ( .D(n178), .CK(clk), .RN(n24), .Q(\gbuff[1][0] )
         );
  DFFRX1 \gbuff_reg[30][31]  ( .D(n1137), .CK(clk), .RN(n18), .Q(
        \gbuff[30][31] ) );
  DFFRX1 \gbuff_reg[30][30]  ( .D(n1136), .CK(clk), .RN(n23), .Q(
        \gbuff[30][30] ) );
  DFFRX1 \gbuff_reg[30][29]  ( .D(n1135), .CK(clk), .RN(n26), .Q(
        \gbuff[30][29] ) );
  DFFRX1 \gbuff_reg[30][28]  ( .D(n1134), .CK(clk), .RN(n18), .Q(
        \gbuff[30][28] ) );
  DFFRX1 \gbuff_reg[30][27]  ( .D(n1133), .CK(clk), .RN(n25), .Q(
        \gbuff[30][27] ) );
  DFFRX1 \gbuff_reg[30][26]  ( .D(n1132), .CK(clk), .RN(n18), .Q(
        \gbuff[30][26] ) );
  DFFRX1 \gbuff_reg[30][25]  ( .D(n1131), .CK(clk), .RN(n24), .Q(
        \gbuff[30][25] ) );
  DFFRX1 \gbuff_reg[30][24]  ( .D(n1130), .CK(clk), .RN(n21), .Q(
        \gbuff[30][24] ) );
  DFFRX1 \gbuff_reg[30][23]  ( .D(n1129), .CK(clk), .RN(n18), .Q(
        \gbuff[30][23] ) );
  DFFRX1 \gbuff_reg[30][22]  ( .D(n1128), .CK(clk), .RN(n23), .Q(
        \gbuff[30][22] ) );
  DFFRX1 \gbuff_reg[30][21]  ( .D(n1127), .CK(clk), .RN(n18), .Q(
        \gbuff[30][21] ) );
  DFFRX1 \gbuff_reg[30][20]  ( .D(n1126), .CK(clk), .RN(n25), .Q(
        \gbuff[30][20] ) );
  DFFRX1 \gbuff_reg[30][19]  ( .D(n1125), .CK(clk), .RN(n17), .Q(
        \gbuff[30][19] ) );
  DFFRX1 \gbuff_reg[30][18]  ( .D(n1124), .CK(clk), .RN(n20), .Q(
        \gbuff[30][18] ) );
  DFFRX1 \gbuff_reg[30][17]  ( .D(n1123), .CK(clk), .RN(n19), .Q(
        \gbuff[30][17] ) );
  DFFRX1 \gbuff_reg[30][16]  ( .D(n1122), .CK(clk), .RN(n17), .Q(
        \gbuff[30][16] ) );
  DFFRX1 \gbuff_reg[30][15]  ( .D(n1121), .CK(clk), .RN(n23), .Q(
        \gbuff[30][15] ) );
  DFFRX1 \gbuff_reg[30][14]  ( .D(n1120), .CK(clk), .RN(n24), .Q(
        \gbuff[30][14] ) );
  DFFRX1 \gbuff_reg[30][13]  ( .D(n1119), .CK(clk), .RN(n24), .Q(
        \gbuff[30][13] ) );
  DFFRX1 \gbuff_reg[30][12]  ( .D(n1118), .CK(clk), .RN(n21), .Q(
        \gbuff[30][12] ) );
  DFFRX1 \gbuff_reg[30][11]  ( .D(n1117), .CK(clk), .RN(n17), .Q(
        \gbuff[30][11] ) );
  DFFRX1 \gbuff_reg[30][10]  ( .D(n1116), .CK(clk), .RN(n24), .Q(
        \gbuff[30][10] ) );
  DFFRX1 \gbuff_reg[30][9]  ( .D(n1115), .CK(clk), .RN(n19), .Q(\gbuff[30][9] ) );
  DFFRX1 \gbuff_reg[30][8]  ( .D(n1114), .CK(clk), .RN(n17), .Q(\gbuff[30][8] ) );
  DFFRX1 \gbuff_reg[30][7]  ( .D(n1113), .CK(clk), .RN(n24), .Q(\gbuff[30][7] ) );
  DFFRX1 \gbuff_reg[30][6]  ( .D(n1112), .CK(clk), .RN(n25), .Q(\gbuff[30][6] ) );
  DFFRX1 \gbuff_reg[30][5]  ( .D(n1111), .CK(clk), .RN(n24), .Q(\gbuff[30][5] ) );
  DFFRX1 \gbuff_reg[30][4]  ( .D(n1110), .CK(clk), .RN(n17), .Q(\gbuff[30][4] ) );
  DFFRX1 \gbuff_reg[30][3]  ( .D(n1109), .CK(clk), .RN(n19), .Q(\gbuff[30][3] ) );
  DFFRX1 \gbuff_reg[30][2]  ( .D(n1108), .CK(clk), .RN(n19), .Q(\gbuff[30][2] ) );
  DFFRX1 \gbuff_reg[30][1]  ( .D(n1107), .CK(clk), .RN(n18), .Q(\gbuff[30][1] ) );
  DFFRX1 \gbuff_reg[30][0]  ( .D(n1106), .CK(clk), .RN(n19), .Q(\gbuff[30][0] ) );
  DFFRX1 \gbuff_reg[26][31]  ( .D(n1009), .CK(clk), .RN(n24), .Q(
        \gbuff[26][31] ) );
  DFFRX1 \gbuff_reg[26][30]  ( .D(n1008), .CK(clk), .RN(n25), .Q(
        \gbuff[26][30] ) );
  DFFRX1 \gbuff_reg[26][29]  ( .D(n1007), .CK(clk), .RN(n20), .Q(
        \gbuff[26][29] ) );
  DFFRX1 \gbuff_reg[26][28]  ( .D(n1006), .CK(clk), .RN(n24), .Q(
        \gbuff[26][28] ) );
  DFFRX1 \gbuff_reg[26][27]  ( .D(n1005), .CK(clk), .RN(n26), .Q(
        \gbuff[26][27] ) );
  DFFRX1 \gbuff_reg[26][26]  ( .D(n1004), .CK(clk), .RN(n23), .Q(
        \gbuff[26][26] ) );
  DFFRX1 \gbuff_reg[26][25]  ( .D(n1003), .CK(clk), .RN(n24), .Q(
        \gbuff[26][25] ) );
  DFFRX1 \gbuff_reg[26][24]  ( .D(n1002), .CK(clk), .RN(n18), .Q(
        \gbuff[26][24] ) );
  DFFRX1 \gbuff_reg[26][23]  ( .D(n1001), .CK(clk), .RN(n21), .Q(
        \gbuff[26][23] ) );
  DFFRX1 \gbuff_reg[26][22]  ( .D(n1000), .CK(clk), .RN(n17), .Q(
        \gbuff[26][22] ) );
  DFFRX1 \gbuff_reg[26][21]  ( .D(n999), .CK(clk), .RN(n17), .Q(
        \gbuff[26][21] ) );
  DFFRX1 \gbuff_reg[26][20]  ( .D(n998), .CK(clk), .RN(n20), .Q(
        \gbuff[26][20] ) );
  DFFRX1 \gbuff_reg[26][19]  ( .D(n997), .CK(clk), .RN(n26), .Q(
        \gbuff[26][19] ) );
  DFFRX1 \gbuff_reg[26][18]  ( .D(n996), .CK(clk), .RN(n26), .Q(
        \gbuff[26][18] ) );
  DFFRX1 \gbuff_reg[26][17]  ( .D(n995), .CK(clk), .RN(n21), .Q(
        \gbuff[26][17] ) );
  DFFRX1 \gbuff_reg[26][16]  ( .D(n994), .CK(clk), .RN(n18), .Q(
        \gbuff[26][16] ) );
  DFFRX1 \gbuff_reg[26][15]  ( .D(n993), .CK(clk), .RN(n25), .Q(
        \gbuff[26][15] ) );
  DFFRX1 \gbuff_reg[26][14]  ( .D(n992), .CK(clk), .RN(n26), .Q(
        \gbuff[26][14] ) );
  DFFRX1 \gbuff_reg[26][13]  ( .D(n991), .CK(clk), .RN(n17), .Q(
        \gbuff[26][13] ) );
  DFFRX1 \gbuff_reg[26][12]  ( .D(n990), .CK(clk), .RN(n20), .Q(
        \gbuff[26][12] ) );
  DFFRX1 \gbuff_reg[26][11]  ( .D(n989), .CK(clk), .RN(n20), .Q(
        \gbuff[26][11] ) );
  DFFRX1 \gbuff_reg[26][10]  ( .D(n988), .CK(clk), .RN(n20), .Q(
        \gbuff[26][10] ) );
  DFFRX1 \gbuff_reg[26][9]  ( .D(n987), .CK(clk), .RN(n17), .Q(\gbuff[26][9] )
         );
  DFFRX1 \gbuff_reg[26][8]  ( .D(n986), .CK(clk), .RN(n23), .Q(\gbuff[26][8] )
         );
  DFFRX1 \gbuff_reg[26][7]  ( .D(n985), .CK(clk), .RN(n25), .Q(\gbuff[26][7] )
         );
  DFFRX1 \gbuff_reg[26][6]  ( .D(n984), .CK(clk), .RN(n26), .Q(\gbuff[26][6] )
         );
  DFFRX1 \gbuff_reg[26][5]  ( .D(n983), .CK(clk), .RN(n21), .Q(\gbuff[26][5] )
         );
  DFFRX1 \gbuff_reg[26][4]  ( .D(n982), .CK(clk), .RN(n26), .Q(\gbuff[26][4] )
         );
  DFFRX1 \gbuff_reg[26][3]  ( .D(n981), .CK(clk), .RN(n23), .Q(\gbuff[26][3] )
         );
  DFFRX1 \gbuff_reg[26][2]  ( .D(n980), .CK(clk), .RN(n21), .Q(\gbuff[26][2] )
         );
  DFFRX1 \gbuff_reg[26][1]  ( .D(n979), .CK(clk), .RN(n23), .Q(\gbuff[26][1] )
         );
  DFFRX1 \gbuff_reg[26][0]  ( .D(n978), .CK(clk), .RN(n20), .Q(\gbuff[26][0] )
         );
  DFFRX1 \gbuff_reg[22][31]  ( .D(n881), .CK(clk), .RN(n18), .Q(
        \gbuff[22][31] ) );
  DFFRX1 \gbuff_reg[22][30]  ( .D(n880), .CK(clk), .RN(n18), .Q(
        \gbuff[22][30] ) );
  DFFRX1 \gbuff_reg[22][29]  ( .D(n879), .CK(clk), .RN(n18), .Q(
        \gbuff[22][29] ) );
  DFFRX1 \gbuff_reg[22][28]  ( .D(n878), .CK(clk), .RN(n18), .Q(
        \gbuff[22][28] ) );
  DFFRX1 \gbuff_reg[22][27]  ( .D(n877), .CK(clk), .RN(n23), .Q(
        \gbuff[22][27] ) );
  DFFRX1 \gbuff_reg[22][26]  ( .D(n876), .CK(clk), .RN(n25), .Q(
        \gbuff[22][26] ) );
  DFFRX1 \gbuff_reg[22][25]  ( .D(n875), .CK(clk), .RN(n20), .Q(
        \gbuff[22][25] ) );
  DFFRX1 \gbuff_reg[22][24]  ( .D(n874), .CK(clk), .RN(n20), .Q(
        \gbuff[22][24] ) );
  DFFRX1 \gbuff_reg[22][23]  ( .D(n873), .CK(clk), .RN(n19), .Q(
        \gbuff[22][23] ) );
  DFFRX1 \gbuff_reg[22][22]  ( .D(n872), .CK(clk), .RN(n24), .Q(
        \gbuff[22][22] ) );
  DFFRX1 \gbuff_reg[22][21]  ( .D(n871), .CK(clk), .RN(n18), .Q(
        \gbuff[22][21] ) );
  DFFRX1 \gbuff_reg[22][20]  ( .D(n870), .CK(clk), .RN(n18), .Q(
        \gbuff[22][20] ) );
  DFFRX1 \gbuff_reg[22][19]  ( .D(n869), .CK(clk), .RN(n17), .Q(
        \gbuff[22][19] ) );
  DFFRX1 \gbuff_reg[22][18]  ( .D(n868), .CK(clk), .RN(n23), .Q(
        \gbuff[22][18] ) );
  DFFRX1 \gbuff_reg[22][17]  ( .D(n867), .CK(clk), .RN(n20), .Q(
        \gbuff[22][17] ) );
  DFFRX1 \gbuff_reg[22][16]  ( .D(n866), .CK(clk), .RN(n25), .Q(
        \gbuff[22][16] ) );
  DFFRX1 \gbuff_reg[22][15]  ( .D(n865), .CK(clk), .RN(n19), .Q(
        \gbuff[22][15] ) );
  DFFRX1 \gbuff_reg[22][14]  ( .D(n864), .CK(clk), .RN(n24), .Q(
        \gbuff[22][14] ) );
  DFFRX1 \gbuff_reg[22][13]  ( .D(n863), .CK(clk), .RN(n19), .Q(
        \gbuff[22][13] ) );
  DFFRX1 \gbuff_reg[22][12]  ( .D(n862), .CK(clk), .RN(n17), .Q(
        \gbuff[22][12] ) );
  DFFRX1 \gbuff_reg[22][11]  ( .D(n861), .CK(clk), .RN(n21), .Q(
        \gbuff[22][11] ) );
  DFFRX1 \gbuff_reg[22][10]  ( .D(n860), .CK(clk), .RN(n25), .Q(
        \gbuff[22][10] ) );
  DFFRX1 \gbuff_reg[22][9]  ( .D(n859), .CK(clk), .RN(n17), .Q(\gbuff[22][9] )
         );
  DFFRX1 \gbuff_reg[22][8]  ( .D(n858), .CK(clk), .RN(n21), .Q(\gbuff[22][8] )
         );
  DFFRX1 \gbuff_reg[22][7]  ( .D(n857), .CK(clk), .RN(n24), .Q(\gbuff[22][7] )
         );
  DFFRX1 \gbuff_reg[22][6]  ( .D(n856), .CK(clk), .RN(n20), .Q(\gbuff[22][6] )
         );
  DFFRX1 \gbuff_reg[22][5]  ( .D(n855), .CK(clk), .RN(n20), .Q(\gbuff[22][5] )
         );
  DFFRX1 \gbuff_reg[22][4]  ( .D(n854), .CK(clk), .RN(n17), .Q(\gbuff[22][4] )
         );
  DFFRX1 \gbuff_reg[22][3]  ( .D(n853), .CK(clk), .RN(n21), .Q(\gbuff[22][3] )
         );
  DFFRX1 \gbuff_reg[22][2]  ( .D(n852), .CK(clk), .RN(n23), .Q(\gbuff[22][2] )
         );
  DFFRX1 \gbuff_reg[22][1]  ( .D(n851), .CK(clk), .RN(n18), .Q(\gbuff[22][1] )
         );
  DFFRX1 \gbuff_reg[22][0]  ( .D(n850), .CK(clk), .RN(n21), .Q(\gbuff[22][0] )
         );
  DFFRX1 \gbuff_reg[18][31]  ( .D(n753), .CK(clk), .RN(n20), .Q(
        \gbuff[18][31] ) );
  DFFRX1 \gbuff_reg[18][30]  ( .D(n752), .CK(clk), .RN(n17), .Q(
        \gbuff[18][30] ) );
  DFFRX1 \gbuff_reg[18][29]  ( .D(n751), .CK(clk), .RN(n20), .Q(
        \gbuff[18][29] ) );
  DFFRX1 \gbuff_reg[18][28]  ( .D(n750), .CK(clk), .RN(n21), .Q(
        \gbuff[18][28] ) );
  DFFRX1 \gbuff_reg[18][27]  ( .D(n749), .CK(clk), .RN(n26), .Q(
        \gbuff[18][27] ) );
  DFFRX1 \gbuff_reg[18][26]  ( .D(n748), .CK(clk), .RN(n21), .Q(
        \gbuff[18][26] ) );
  DFFRX1 \gbuff_reg[18][25]  ( .D(n747), .CK(clk), .RN(n18), .Q(
        \gbuff[18][25] ) );
  DFFRX1 \gbuff_reg[18][24]  ( .D(n746), .CK(clk), .RN(n26), .Q(
        \gbuff[18][24] ) );
  DFFRX1 \gbuff_reg[18][23]  ( .D(n745), .CK(clk), .RN(n20), .Q(
        \gbuff[18][23] ) );
  DFFRX1 \gbuff_reg[18][22]  ( .D(n744), .CK(clk), .RN(n17), .Q(
        \gbuff[18][22] ) );
  DFFRX1 \gbuff_reg[18][21]  ( .D(n743), .CK(clk), .RN(n23), .Q(
        \gbuff[18][21] ) );
  DFFRX1 \gbuff_reg[18][20]  ( .D(n742), .CK(clk), .RN(n24), .Q(
        \gbuff[18][20] ) );
  DFFRX1 \gbuff_reg[18][19]  ( .D(n741), .CK(clk), .RN(n18), .Q(
        \gbuff[18][19] ) );
  DFFRX1 \gbuff_reg[18][18]  ( .D(n740), .CK(clk), .RN(n19), .Q(
        \gbuff[18][18] ) );
  DFFRX1 \gbuff_reg[18][17]  ( .D(n739), .CK(clk), .RN(n25), .Q(
        \gbuff[18][17] ) );
  DFFRX1 \gbuff_reg[18][16]  ( .D(n738), .CK(clk), .RN(n19), .Q(
        \gbuff[18][16] ) );
  DFFRX1 \gbuff_reg[18][15]  ( .D(n737), .CK(clk), .RN(n25), .Q(
        \gbuff[18][15] ) );
  DFFRX1 \gbuff_reg[18][14]  ( .D(n736), .CK(clk), .RN(n21), .Q(
        \gbuff[18][14] ) );
  DFFRX1 \gbuff_reg[18][13]  ( .D(n735), .CK(clk), .RN(n21), .Q(
        \gbuff[18][13] ) );
  DFFRX1 \gbuff_reg[18][12]  ( .D(n734), .CK(clk), .RN(n24), .Q(
        \gbuff[18][12] ) );
  DFFRX1 \gbuff_reg[18][11]  ( .D(n733), .CK(clk), .RN(n18), .Q(
        \gbuff[18][11] ) );
  DFFRX1 \gbuff_reg[18][10]  ( .D(n732), .CK(clk), .RN(n19), .Q(
        \gbuff[18][10] ) );
  DFFRX1 \gbuff_reg[18][9]  ( .D(n731), .CK(clk), .RN(n17), .Q(\gbuff[18][9] )
         );
  DFFRX1 \gbuff_reg[18][8]  ( .D(n730), .CK(clk), .RN(n19), .Q(\gbuff[18][8] )
         );
  DFFRX1 \gbuff_reg[18][7]  ( .D(n729), .CK(clk), .RN(n17), .Q(\gbuff[18][7] )
         );
  DFFRX1 \gbuff_reg[18][6]  ( .D(n728), .CK(clk), .RN(n18), .Q(\gbuff[18][6] )
         );
  DFFRX1 \gbuff_reg[18][5]  ( .D(n727), .CK(clk), .RN(n21), .Q(\gbuff[18][5] )
         );
  DFFRX1 \gbuff_reg[18][4]  ( .D(n726), .CK(clk), .RN(n20), .Q(\gbuff[18][4] )
         );
  DFFRX1 \gbuff_reg[18][3]  ( .D(n725), .CK(clk), .RN(n23), .Q(\gbuff[18][3] )
         );
  DFFRX1 \gbuff_reg[18][2]  ( .D(n724), .CK(clk), .RN(n25), .Q(\gbuff[18][2] )
         );
  DFFRX1 \gbuff_reg[18][1]  ( .D(n723), .CK(clk), .RN(n21), .Q(\gbuff[18][1] )
         );
  DFFRX1 \gbuff_reg[18][0]  ( .D(n722), .CK(clk), .RN(n24), .Q(\gbuff[18][0] )
         );
  DFFRX1 \gbuff_reg[14][31]  ( .D(n625), .CK(clk), .RN(n17), .Q(
        \gbuff[14][31] ) );
  DFFRX1 \gbuff_reg[14][30]  ( .D(n624), .CK(clk), .RN(n18), .Q(
        \gbuff[14][30] ) );
  DFFRX1 \gbuff_reg[14][29]  ( .D(n623), .CK(clk), .RN(n25), .Q(
        \gbuff[14][29] ) );
  DFFRX1 \gbuff_reg[14][28]  ( .D(n622), .CK(clk), .RN(n18), .Q(
        \gbuff[14][28] ) );
  DFFRX1 \gbuff_reg[14][27]  ( .D(n621), .CK(clk), .RN(n24), .Q(
        \gbuff[14][27] ) );
  DFFRX1 \gbuff_reg[14][26]  ( .D(n620), .CK(clk), .RN(n26), .Q(
        \gbuff[14][26] ) );
  DFFRX1 \gbuff_reg[14][25]  ( .D(n619), .CK(clk), .RN(n18), .Q(
        \gbuff[14][25] ) );
  DFFRX1 \gbuff_reg[14][24]  ( .D(n618), .CK(clk), .RN(n23), .Q(
        \gbuff[14][24] ) );
  DFFRX1 \gbuff_reg[14][23]  ( .D(n617), .CK(clk), .RN(n19), .Q(
        \gbuff[14][23] ) );
  DFFRX1 \gbuff_reg[14][22]  ( .D(n616), .CK(clk), .RN(n19), .Q(
        \gbuff[14][22] ) );
  DFFRX1 \gbuff_reg[14][21]  ( .D(n615), .CK(clk), .RN(n19), .Q(
        \gbuff[14][21] ) );
  DFFRX1 \gbuff_reg[14][20]  ( .D(n614), .CK(clk), .RN(n26), .Q(
        \gbuff[14][20] ) );
  DFFRX1 \gbuff_reg[14][19]  ( .D(n613), .CK(clk), .RN(n24), .Q(
        \gbuff[14][19] ) );
  DFFRX1 \gbuff_reg[14][18]  ( .D(n612), .CK(clk), .RN(n21), .Q(
        \gbuff[14][18] ) );
  DFFRX1 \gbuff_reg[14][17]  ( .D(n611), .CK(clk), .RN(n24), .Q(
        \gbuff[14][17] ) );
  DFFRX1 \gbuff_reg[14][16]  ( .D(n610), .CK(clk), .RN(n23), .Q(
        \gbuff[14][16] ) );
  DFFRX1 \gbuff_reg[14][15]  ( .D(n609), .CK(clk), .RN(n26), .Q(
        \gbuff[14][15] ) );
  DFFRX1 \gbuff_reg[14][14]  ( .D(n608), .CK(clk), .RN(n20), .Q(
        \gbuff[14][14] ) );
  DFFRX1 \gbuff_reg[14][13]  ( .D(n607), .CK(clk), .RN(n19), .Q(
        \gbuff[14][13] ) );
  DFFRX1 \gbuff_reg[14][12]  ( .D(n606), .CK(clk), .RN(n19), .Q(
        \gbuff[14][12] ) );
  DFFRX1 \gbuff_reg[14][11]  ( .D(n605), .CK(clk), .RN(n21), .Q(
        \gbuff[14][11] ) );
  DFFRX1 \gbuff_reg[14][10]  ( .D(n604), .CK(clk), .RN(n19), .Q(
        \gbuff[14][10] ) );
  DFFRX1 \gbuff_reg[14][9]  ( .D(n603), .CK(clk), .RN(n20), .Q(\gbuff[14][9] )
         );
  DFFRX1 \gbuff_reg[14][8]  ( .D(n602), .CK(clk), .RN(n17), .Q(\gbuff[14][8] )
         );
  DFFRX1 \gbuff_reg[14][7]  ( .D(n601), .CK(clk), .RN(n26), .Q(\gbuff[14][7] )
         );
  DFFRX1 \gbuff_reg[14][6]  ( .D(n600), .CK(clk), .RN(n20), .Q(\gbuff[14][6] )
         );
  DFFRX1 \gbuff_reg[14][5]  ( .D(n599), .CK(clk), .RN(n26), .Q(\gbuff[14][5] )
         );
  DFFRX1 \gbuff_reg[14][4]  ( .D(n598), .CK(clk), .RN(n17), .Q(\gbuff[14][4] )
         );
  DFFRX1 \gbuff_reg[14][3]  ( .D(n597), .CK(clk), .RN(n25), .Q(\gbuff[14][3] )
         );
  DFFRX1 \gbuff_reg[14][2]  ( .D(n596), .CK(clk), .RN(n23), .Q(\gbuff[14][2] )
         );
  DFFRX1 \gbuff_reg[14][1]  ( .D(n595), .CK(clk), .RN(n26), .Q(\gbuff[14][1] )
         );
  DFFRX1 \gbuff_reg[14][0]  ( .D(n594), .CK(clk), .RN(n25), .Q(\gbuff[14][0] )
         );
  DFFRX1 \gbuff_reg[10][31]  ( .D(n497), .CK(clk), .RN(n20), .Q(
        \gbuff[10][31] ) );
  DFFRX1 \gbuff_reg[10][30]  ( .D(n496), .CK(clk), .RN(n23), .Q(
        \gbuff[10][30] ) );
  DFFRX1 \gbuff_reg[10][29]  ( .D(n495), .CK(clk), .RN(n23), .Q(
        \gbuff[10][29] ) );
  DFFRX1 \gbuff_reg[10][28]  ( .D(n494), .CK(clk), .RN(n25), .Q(
        \gbuff[10][28] ) );
  DFFRX1 \gbuff_reg[10][27]  ( .D(n493), .CK(clk), .RN(n25), .Q(
        \gbuff[10][27] ) );
  DFFRX1 \gbuff_reg[10][26]  ( .D(n492), .CK(clk), .RN(n20), .Q(
        \gbuff[10][26] ) );
  DFFRX1 \gbuff_reg[10][25]  ( .D(n491), .CK(clk), .RN(n26), .Q(
        \gbuff[10][25] ) );
  DFFRX1 \gbuff_reg[10][24]  ( .D(n490), .CK(clk), .RN(n25), .Q(
        \gbuff[10][24] ) );
  DFFRX1 \gbuff_reg[10][23]  ( .D(n489), .CK(clk), .RN(n23), .Q(
        \gbuff[10][23] ) );
  DFFRX1 \gbuff_reg[10][22]  ( .D(n488), .CK(clk), .RN(n21), .Q(
        \gbuff[10][22] ) );
  DFFRX1 \gbuff_reg[10][21]  ( .D(n487), .CK(clk), .RN(n23), .Q(
        \gbuff[10][21] ) );
  DFFRX1 \gbuff_reg[10][20]  ( .D(n486), .CK(clk), .RN(n21), .Q(
        \gbuff[10][20] ) );
  DFFRX1 \gbuff_reg[10][19]  ( .D(n485), .CK(clk), .RN(n18), .Q(
        \gbuff[10][19] ) );
  DFFRX1 \gbuff_reg[10][18]  ( .D(n484), .CK(clk), .RN(n26), .Q(
        \gbuff[10][18] ) );
  DFFRX1 \gbuff_reg[10][17]  ( .D(n483), .CK(clk), .RN(n19), .Q(
        \gbuff[10][17] ) );
  DFFRX1 \gbuff_reg[10][16]  ( .D(n482), .CK(clk), .RN(n18), .Q(
        \gbuff[10][16] ) );
  DFFRX1 \gbuff_reg[10][15]  ( .D(n481), .CK(clk), .RN(n23), .Q(
        \gbuff[10][15] ) );
  DFFRX1 \gbuff_reg[10][14]  ( .D(n480), .CK(clk), .RN(n21), .Q(
        \gbuff[10][14] ) );
  DFFRX1 \gbuff_reg[10][13]  ( .D(n479), .CK(clk), .RN(n24), .Q(
        \gbuff[10][13] ) );
  DFFRX1 \gbuff_reg[10][12]  ( .D(n478), .CK(clk), .RN(n20), .Q(
        \gbuff[10][12] ) );
  DFFRX1 \gbuff_reg[10][11]  ( .D(n477), .CK(clk), .RN(n19), .Q(
        \gbuff[10][11] ) );
  DFFRX1 \gbuff_reg[10][10]  ( .D(n476), .CK(clk), .RN(n24), .Q(
        \gbuff[10][10] ) );
  DFFRX1 \gbuff_reg[10][9]  ( .D(n475), .CK(clk), .RN(n20), .Q(\gbuff[10][9] )
         );
  DFFRX1 \gbuff_reg[10][8]  ( .D(n474), .CK(clk), .RN(n26), .Q(\gbuff[10][8] )
         );
  DFFRX1 \gbuff_reg[10][7]  ( .D(n473), .CK(clk), .RN(n17), .Q(\gbuff[10][7] )
         );
  DFFRX1 \gbuff_reg[10][6]  ( .D(n472), .CK(clk), .RN(n25), .Q(\gbuff[10][6] )
         );
  DFFRX1 \gbuff_reg[10][5]  ( .D(n471), .CK(clk), .RN(n25), .Q(\gbuff[10][5] )
         );
  DFFRX1 \gbuff_reg[10][4]  ( .D(n470), .CK(clk), .RN(n23), .Q(\gbuff[10][4] )
         );
  DFFRX1 \gbuff_reg[10][3]  ( .D(n469), .CK(clk), .RN(n19), .Q(\gbuff[10][3] )
         );
  DFFRX1 \gbuff_reg[10][2]  ( .D(n468), .CK(clk), .RN(n18), .Q(\gbuff[10][2] )
         );
  DFFRX1 \gbuff_reg[10][1]  ( .D(n467), .CK(clk), .RN(n25), .Q(\gbuff[10][1] )
         );
  DFFRX1 \gbuff_reg[10][0]  ( .D(n466), .CK(clk), .RN(n26), .Q(\gbuff[10][0] )
         );
  DFFRX1 \gbuff_reg[6][31]  ( .D(n369), .CK(clk), .RN(n21), .Q(\gbuff[6][31] )
         );
  DFFRX1 \gbuff_reg[6][30]  ( .D(n368), .CK(clk), .RN(n19), .Q(\gbuff[6][30] )
         );
  DFFRX1 \gbuff_reg[6][29]  ( .D(n367), .CK(clk), .RN(n25), .Q(\gbuff[6][29] )
         );
  DFFRX1 \gbuff_reg[6][28]  ( .D(n366), .CK(clk), .RN(n23), .Q(\gbuff[6][28] )
         );
  DFFRX1 \gbuff_reg[6][27]  ( .D(n365), .CK(clk), .RN(n24), .Q(\gbuff[6][27] )
         );
  DFFRX1 \gbuff_reg[6][26]  ( .D(n364), .CK(clk), .RN(n23), .Q(\gbuff[6][26] )
         );
  DFFRX1 \gbuff_reg[6][25]  ( .D(n363), .CK(clk), .RN(n21), .Q(\gbuff[6][25] )
         );
  DFFRX1 \gbuff_reg[6][24]  ( .D(n362), .CK(clk), .RN(n20), .Q(\gbuff[6][24] )
         );
  DFFRX1 \gbuff_reg[6][23]  ( .D(n361), .CK(clk), .RN(n21), .Q(\gbuff[6][23] )
         );
  DFFRX1 \gbuff_reg[6][22]  ( .D(n360), .CK(clk), .RN(n19), .Q(\gbuff[6][22] )
         );
  DFFRX1 \gbuff_reg[6][21]  ( .D(n359), .CK(clk), .RN(n17), .Q(\gbuff[6][21] )
         );
  DFFRX1 \gbuff_reg[6][20]  ( .D(n358), .CK(clk), .RN(n18), .Q(\gbuff[6][20] )
         );
  DFFRX1 \gbuff_reg[6][19]  ( .D(n357), .CK(clk), .RN(n20), .Q(\gbuff[6][19] )
         );
  DFFRX1 \gbuff_reg[6][18]  ( .D(n356), .CK(clk), .RN(n25), .Q(\gbuff[6][18] )
         );
  DFFRX1 \gbuff_reg[6][17]  ( .D(n355), .CK(clk), .RN(n24), .Q(\gbuff[6][17] )
         );
  DFFRX1 \gbuff_reg[6][16]  ( .D(n354), .CK(clk), .RN(n24), .Q(\gbuff[6][16] )
         );
  DFFRX1 \gbuff_reg[6][15]  ( .D(n353), .CK(clk), .RN(n26), .Q(\gbuff[6][15] )
         );
  DFFRX1 \gbuff_reg[6][14]  ( .D(n352), .CK(clk), .RN(n26), .Q(\gbuff[6][14] )
         );
  DFFRX1 \gbuff_reg[6][13]  ( .D(n351), .CK(clk), .RN(n26), .Q(\gbuff[6][13] )
         );
  DFFRX1 \gbuff_reg[6][12]  ( .D(n350), .CK(clk), .RN(n19), .Q(\gbuff[6][12] )
         );
  DFFRX1 \gbuff_reg[6][11]  ( .D(n349), .CK(clk), .RN(n20), .Q(\gbuff[6][11] )
         );
  DFFRX1 \gbuff_reg[6][10]  ( .D(n348), .CK(clk), .RN(n17), .Q(\gbuff[6][10] )
         );
  DFFRX1 \gbuff_reg[6][9]  ( .D(n347), .CK(clk), .RN(n23), .Q(\gbuff[6][9] )
         );
  DFFRX1 \gbuff_reg[6][8]  ( .D(n346), .CK(clk), .RN(n24), .Q(\gbuff[6][8] )
         );
  DFFRX1 \gbuff_reg[6][7]  ( .D(n345), .CK(clk), .RN(n18), .Q(\gbuff[6][7] )
         );
  DFFRX1 \gbuff_reg[6][6]  ( .D(n344), .CK(clk), .RN(n23), .Q(\gbuff[6][6] )
         );
  DFFRX1 \gbuff_reg[6][5]  ( .D(n343), .CK(clk), .RN(n26), .Q(\gbuff[6][5] )
         );
  DFFRX1 \gbuff_reg[6][4]  ( .D(n342), .CK(clk), .RN(n19), .Q(\gbuff[6][4] )
         );
  DFFRX1 \gbuff_reg[6][3]  ( .D(n341), .CK(clk), .RN(n25), .Q(\gbuff[6][3] )
         );
  DFFRX1 \gbuff_reg[6][2]  ( .D(n340), .CK(clk), .RN(n24), .Q(\gbuff[6][2] )
         );
  DFFRX1 \gbuff_reg[6][1]  ( .D(n339), .CK(clk), .RN(n23), .Q(\gbuff[6][1] )
         );
  DFFRX1 \gbuff_reg[6][0]  ( .D(n338), .CK(clk), .RN(n21), .Q(\gbuff[6][0] )
         );
  DFFRX1 \gbuff_reg[2][31]  ( .D(n241), .CK(clk), .RN(n18), .Q(\gbuff[2][31] )
         );
  DFFRX1 \gbuff_reg[2][30]  ( .D(n240), .CK(clk), .RN(n23), .Q(\gbuff[2][30] )
         );
  DFFRX1 \gbuff_reg[2][29]  ( .D(n239), .CK(clk), .RN(n18), .Q(\gbuff[2][29] )
         );
  DFFRX1 \gbuff_reg[2][28]  ( .D(n238), .CK(clk), .RN(n21), .Q(\gbuff[2][28] )
         );
  DFFRX1 \gbuff_reg[2][27]  ( .D(n237), .CK(clk), .RN(n17), .Q(\gbuff[2][27] )
         );
  DFFRX1 \gbuff_reg[2][26]  ( .D(n236), .CK(clk), .RN(n17), .Q(\gbuff[2][26] )
         );
  DFFRX1 \gbuff_reg[2][25]  ( .D(n235), .CK(clk), .RN(n21), .Q(\gbuff[2][25] )
         );
  DFFRX1 \gbuff_reg[2][24]  ( .D(n234), .CK(clk), .RN(n17), .Q(\gbuff[2][24] )
         );
  DFFRX1 \gbuff_reg[2][23]  ( .D(n233), .CK(clk), .RN(n23), .Q(\gbuff[2][23] )
         );
  DFFRX1 \gbuff_reg[2][22]  ( .D(n232), .CK(clk), .RN(n24), .Q(\gbuff[2][22] )
         );
  DFFRX1 \gbuff_reg[2][21]  ( .D(n231), .CK(clk), .RN(n24), .Q(\gbuff[2][21] )
         );
  DFFRX1 \gbuff_reg[2][20]  ( .D(n230), .CK(clk), .RN(n21), .Q(\gbuff[2][20] )
         );
  DFFRX1 \gbuff_reg[2][19]  ( .D(n229), .CK(clk), .RN(n17), .Q(\gbuff[2][19] )
         );
  DFFRX1 \gbuff_reg[2][18]  ( .D(n228), .CK(clk), .RN(n24), .Q(\gbuff[2][18] )
         );
  DFFRX1 \gbuff_reg[2][17]  ( .D(n227), .CK(clk), .RN(n19), .Q(\gbuff[2][17] )
         );
  DFFRX1 \gbuff_reg[2][16]  ( .D(n226), .CK(clk), .RN(n17), .Q(\gbuff[2][16] )
         );
  DFFRX1 \gbuff_reg[2][15]  ( .D(n225), .CK(clk), .RN(n24), .Q(\gbuff[2][15] )
         );
  DFFRX1 \gbuff_reg[2][14]  ( .D(n224), .CK(clk), .RN(n25), .Q(\gbuff[2][14] )
         );
  DFFRX1 \gbuff_reg[2][13]  ( .D(n223), .CK(clk), .RN(n24), .Q(\gbuff[2][13] )
         );
  DFFRX1 \gbuff_reg[2][12]  ( .D(n222), .CK(clk), .RN(n25), .Q(\gbuff[2][12] )
         );
  DFFRX1 \gbuff_reg[2][11]  ( .D(n221), .CK(clk), .RN(n19), .Q(\gbuff[2][11] )
         );
  DFFRX1 \gbuff_reg[2][10]  ( .D(n220), .CK(clk), .RN(n25), .Q(\gbuff[2][10] )
         );
  DFFRX1 \gbuff_reg[2][9]  ( .D(n219), .CK(clk), .RN(n19), .Q(\gbuff[2][9] )
         );
  DFFRX1 \gbuff_reg[2][8]  ( .D(n218), .CK(clk), .RN(n19), .Q(\gbuff[2][8] )
         );
  DFFRX1 \gbuff_reg[2][7]  ( .D(n217), .CK(clk), .RN(n24), .Q(\gbuff[2][7] )
         );
  DFFRX1 \gbuff_reg[2][6]  ( .D(n216), .CK(clk), .RN(n25), .Q(\gbuff[2][6] )
         );
  DFFRX1 \gbuff_reg[2][5]  ( .D(n215), .CK(clk), .RN(n20), .Q(\gbuff[2][5] )
         );
  DFFRX1 \gbuff_reg[2][4]  ( .D(n214), .CK(clk), .RN(n20), .Q(\gbuff[2][4] )
         );
  DFFRX1 \gbuff_reg[2][3]  ( .D(n213), .CK(clk), .RN(n26), .Q(\gbuff[2][3] )
         );
  DFFRX1 \gbuff_reg[2][2]  ( .D(n212), .CK(clk), .RN(n26), .Q(\gbuff[2][2] )
         );
  DFFRX1 \gbuff_reg[2][1]  ( .D(n211), .CK(clk), .RN(n17), .Q(\gbuff[2][1] )
         );
  DFFRX1 \gbuff_reg[2][0]  ( .D(n210), .CK(clk), .RN(n18), .Q(\gbuff[2][0] )
         );
  DFFRX1 \gbuff_reg[28][31]  ( .D(n1073), .CK(clk), .RN(n21), .Q(
        \gbuff[28][31] ) );
  DFFRX1 \gbuff_reg[28][30]  ( .D(n1072), .CK(clk), .RN(n17), .Q(
        \gbuff[28][30] ) );
  DFFRX1 \gbuff_reg[28][29]  ( .D(n1071), .CK(clk), .RN(n17), .Q(
        \gbuff[28][29] ) );
  DFFRX1 \gbuff_reg[28][28]  ( .D(n1070), .CK(clk), .RN(n20), .Q(
        \gbuff[28][28] ) );
  DFFRX1 \gbuff_reg[28][27]  ( .D(n1069), .CK(clk), .RN(n26), .Q(
        \gbuff[28][27] ) );
  DFFRX1 \gbuff_reg[28][26]  ( .D(n1068), .CK(clk), .RN(n26), .Q(
        \gbuff[28][26] ) );
  DFFRX1 \gbuff_reg[28][25]  ( .D(n1067), .CK(clk), .RN(n21), .Q(
        \gbuff[28][25] ) );
  DFFRX1 \gbuff_reg[28][24]  ( .D(n1066), .CK(clk), .RN(n18), .Q(
        \gbuff[28][24] ) );
  DFFRX1 \gbuff_reg[28][23]  ( .D(n1065), .CK(clk), .RN(n25), .Q(
        \gbuff[28][23] ) );
  DFFRX1 \gbuff_reg[28][22]  ( .D(n1064), .CK(clk), .RN(n26), .Q(
        \gbuff[28][22] ) );
  DFFRX1 \gbuff_reg[28][21]  ( .D(n1063), .CK(clk), .RN(n17), .Q(
        \gbuff[28][21] ) );
  DFFRX1 \gbuff_reg[28][20]  ( .D(n1062), .CK(clk), .RN(n23), .Q(
        \gbuff[28][20] ) );
  DFFRX1 \gbuff_reg[28][19]  ( .D(n1061), .CK(clk), .RN(n20), .Q(
        \gbuff[28][19] ) );
  DFFRX1 \gbuff_reg[28][18]  ( .D(n1060), .CK(clk), .RN(n17), .Q(
        \gbuff[28][18] ) );
  DFFRX1 \gbuff_reg[28][17]  ( .D(n1059), .CK(clk), .RN(n25), .Q(
        \gbuff[28][17] ) );
  DFFRX1 \gbuff_reg[28][16]  ( .D(n1058), .CK(clk), .RN(n23), .Q(
        \gbuff[28][16] ) );
  DFFRX1 \gbuff_reg[28][15]  ( .D(n1057), .CK(clk), .RN(n25), .Q(
        \gbuff[28][15] ) );
  DFFRX1 \gbuff_reg[28][14]  ( .D(n1056), .CK(clk), .RN(n26), .Q(
        \gbuff[28][14] ) );
  DFFRX1 \gbuff_reg[28][13]  ( .D(n1055), .CK(clk), .RN(n21), .Q(
        \gbuff[28][13] ) );
  DFFRX1 \gbuff_reg[28][12]  ( .D(n1054), .CK(clk), .RN(n19), .Q(
        \gbuff[28][12] ) );
  DFFRX1 \gbuff_reg[28][11]  ( .D(n1053), .CK(clk), .RN(n23), .Q(
        \gbuff[28][11] ) );
  DFFRX1 \gbuff_reg[28][10]  ( .D(n1052), .CK(clk), .RN(n18), .Q(
        \gbuff[28][10] ) );
  DFFRX1 \gbuff_reg[28][9]  ( .D(n1051), .CK(clk), .RN(n19), .Q(\gbuff[28][9] ) );
  DFFRX1 \gbuff_reg[28][8]  ( .D(n1050), .CK(clk), .RN(n20), .Q(\gbuff[28][8] ) );
  DFFRX1 \gbuff_reg[28][7]  ( .D(n1049), .CK(clk), .RN(n18), .Q(\gbuff[28][7] ) );
  DFFRX1 \gbuff_reg[28][6]  ( .D(n1048), .CK(clk), .RN(n18), .Q(\gbuff[28][6] ) );
  DFFRX1 \gbuff_reg[28][5]  ( .D(n1047), .CK(clk), .RN(n18), .Q(\gbuff[28][5] ) );
  DFFRX1 \gbuff_reg[28][4]  ( .D(n1046), .CK(clk), .RN(n18), .Q(\gbuff[28][4] ) );
  DFFRX1 \gbuff_reg[28][3]  ( .D(n1045), .CK(clk), .RN(n23), .Q(\gbuff[28][3] ) );
  DFFRX1 \gbuff_reg[28][2]  ( .D(n1044), .CK(clk), .RN(n25), .Q(\gbuff[28][2] ) );
  DFFRX1 \gbuff_reg[28][1]  ( .D(n1043), .CK(clk), .RN(n20), .Q(\gbuff[28][1] ) );
  DFFRX1 \gbuff_reg[28][0]  ( .D(n1042), .CK(clk), .RN(n20), .Q(\gbuff[28][0] ) );
  DFFRX1 \gbuff_reg[24][31]  ( .D(n945), .CK(clk), .RN(n19), .Q(
        \gbuff[24][31] ) );
  DFFRX1 \gbuff_reg[24][30]  ( .D(n944), .CK(clk), .RN(n24), .Q(
        \gbuff[24][30] ) );
  DFFRX1 \gbuff_reg[24][29]  ( .D(n943), .CK(clk), .RN(n18), .Q(
        \gbuff[24][29] ) );
  DFFRX1 \gbuff_reg[24][28]  ( .D(n942), .CK(clk), .RN(n26), .Q(
        \gbuff[24][28] ) );
  DFFRX1 \gbuff_reg[24][27]  ( .D(n941), .CK(clk), .RN(n17), .Q(
        \gbuff[24][27] ) );
  DFFRX1 \gbuff_reg[24][26]  ( .D(n940), .CK(clk), .RN(n26), .Q(
        \gbuff[24][26] ) );
  DFFRX1 \gbuff_reg[24][25]  ( .D(n939), .CK(clk), .RN(n23), .Q(
        \gbuff[24][25] ) );
  DFFRX1 \gbuff_reg[24][24]  ( .D(n938), .CK(clk), .RN(n25), .Q(
        \gbuff[24][24] ) );
  DFFRX1 \gbuff_reg[24][23]  ( .D(n937), .CK(clk), .RN(n19), .Q(
        \gbuff[24][23] ) );
  DFFRX1 \gbuff_reg[24][22]  ( .D(n936), .CK(clk), .RN(n24), .Q(
        \gbuff[24][22] ) );
  DFFRX1 \gbuff_reg[24][21]  ( .D(n935), .CK(clk), .RN(n19), .Q(
        \gbuff[24][21] ) );
  DFFRX1 \gbuff_reg[24][20]  ( .D(n934), .CK(clk), .RN(n21), .Q(
        \gbuff[24][20] ) );
  DFFRX1 \gbuff_reg[24][19]  ( .D(n933), .CK(clk), .RN(n21), .Q(
        \gbuff[24][19] ) );
  DFFRX1 \gbuff_reg[24][18]  ( .D(n932), .CK(clk), .RN(n24), .Q(
        \gbuff[24][18] ) );
  DFFRX1 \gbuff_reg[24][17]  ( .D(n931), .CK(clk), .RN(n18), .Q(
        \gbuff[24][17] ) );
  DFFRX1 \gbuff_reg[24][16]  ( .D(n930), .CK(clk), .RN(n21), .Q(
        \gbuff[24][16] ) );
  DFFRX1 \gbuff_reg[24][15]  ( .D(n929), .CK(clk), .RN(n24), .Q(
        \gbuff[24][15] ) );
  DFFRX1 \gbuff_reg[24][14]  ( .D(n928), .CK(clk), .RN(n20), .Q(
        \gbuff[24][14] ) );
  DFFRX1 \gbuff_reg[24][13]  ( .D(n927), .CK(clk), .RN(n20), .Q(
        \gbuff[24][13] ) );
  DFFRX1 \gbuff_reg[24][12]  ( .D(n926), .CK(clk), .RN(n17), .Q(
        \gbuff[24][12] ) );
  DFFRX1 \gbuff_reg[24][11]  ( .D(n925), .CK(clk), .RN(n21), .Q(
        \gbuff[24][11] ) );
  DFFRX1 \gbuff_reg[24][10]  ( .D(n924), .CK(clk), .RN(n23), .Q(
        \gbuff[24][10] ) );
  DFFRX1 \gbuff_reg[24][9]  ( .D(n923), .CK(clk), .RN(n18), .Q(\gbuff[24][9] )
         );
  DFFRX1 \gbuff_reg[24][8]  ( .D(n922), .CK(clk), .RN(n21), .Q(\gbuff[24][8] )
         );
  DFFRX1 \gbuff_reg[24][7]  ( .D(n921), .CK(clk), .RN(n20), .Q(\gbuff[24][7] )
         );
  DFFRX1 \gbuff_reg[24][6]  ( .D(n920), .CK(clk), .RN(n17), .Q(\gbuff[24][6] )
         );
  DFFRX1 \gbuff_reg[24][5]  ( .D(n919), .CK(clk), .RN(n20), .Q(\gbuff[24][5] )
         );
  DFFRX1 \gbuff_reg[24][4]  ( .D(n918), .CK(clk), .RN(n25), .Q(\gbuff[24][4] )
         );
  DFFRX1 \gbuff_reg[24][3]  ( .D(n917), .CK(clk), .RN(n26), .Q(\gbuff[24][3] )
         );
  DFFRX1 \gbuff_reg[24][2]  ( .D(n916), .CK(clk), .RN(n18), .Q(\gbuff[24][2] )
         );
  DFFRX1 \gbuff_reg[24][1]  ( .D(n915), .CK(clk), .RN(n26), .Q(\gbuff[24][1] )
         );
  DFFRX1 \gbuff_reg[24][0]  ( .D(n914), .CK(clk), .RN(n26), .Q(\gbuff[24][0] )
         );
  DFFRX1 \gbuff_reg[20][31]  ( .D(n817), .CK(clk), .RN(n20), .Q(
        \gbuff[20][31] ) );
  DFFRX1 \gbuff_reg[20][30]  ( .D(n816), .CK(clk), .RN(n17), .Q(
        \gbuff[20][30] ) );
  DFFRX1 \gbuff_reg[20][29]  ( .D(n815), .CK(clk), .RN(n23), .Q(
        \gbuff[20][29] ) );
  DFFRX1 \gbuff_reg[20][28]  ( .D(n814), .CK(clk), .RN(n23), .Q(
        \gbuff[20][28] ) );
  DFFRX1 \gbuff_reg[20][27]  ( .D(n813), .CK(clk), .RN(n18), .Q(
        \gbuff[20][27] ) );
  DFFRX1 \gbuff_reg[20][26]  ( .D(n812), .CK(clk), .RN(n20), .Q(
        \gbuff[20][26] ) );
  DFFRX1 \gbuff_reg[20][25]  ( .D(n811), .CK(clk), .RN(n23), .Q(
        \gbuff[20][25] ) );
  DFFRX1 \gbuff_reg[20][24]  ( .D(n810), .CK(clk), .RN(n19), .Q(
        \gbuff[20][24] ) );
  DFFRX1 \gbuff_reg[20][23]  ( .D(n809), .CK(clk), .RN(n25), .Q(
        \gbuff[20][23] ) );
  DFFRX1 \gbuff_reg[20][22]  ( .D(n808), .CK(clk), .RN(n21), .Q(
        \gbuff[20][22] ) );
  DFFRX1 \gbuff_reg[20][21]  ( .D(n807), .CK(clk), .RN(n21), .Q(
        \gbuff[20][21] ) );
  DFFRX1 \gbuff_reg[20][20]  ( .D(n806), .CK(clk), .RN(n24), .Q(
        \gbuff[20][20] ) );
  DFFRX1 \gbuff_reg[20][19]  ( .D(n805), .CK(clk), .RN(n18), .Q(
        \gbuff[20][19] ) );
  DFFRX1 \gbuff_reg[20][18]  ( .D(n804), .CK(clk), .RN(n19), .Q(
        \gbuff[20][18] ) );
  DFFRX1 \gbuff_reg[20][17]  ( .D(n803), .CK(clk), .RN(n17), .Q(
        \gbuff[20][17] ) );
  DFFRX1 \gbuff_reg[20][16]  ( .D(n802), .CK(clk), .RN(n19), .Q(
        \gbuff[20][16] ) );
  DFFRX1 \gbuff_reg[20][15]  ( .D(n801), .CK(clk), .RN(n17), .Q(
        \gbuff[20][15] ) );
  DFFRX1 \gbuff_reg[20][14]  ( .D(n800), .CK(clk), .RN(n18), .Q(
        \gbuff[20][14] ) );
  DFFRX1 \gbuff_reg[20][13]  ( .D(n799), .CK(clk), .RN(n21), .Q(
        \gbuff[20][13] ) );
  DFFRX1 \gbuff_reg[20][12]  ( .D(n798), .CK(clk), .RN(n24), .Q(
        \gbuff[20][12] ) );
  DFFRX1 \gbuff_reg[20][11]  ( .D(n797), .CK(clk), .RN(n23), .Q(
        \gbuff[20][11] ) );
  DFFRX1 \gbuff_reg[20][10]  ( .D(n796), .CK(clk), .RN(n24), .Q(
        \gbuff[20][10] ) );
  DFFRX1 \gbuff_reg[20][9]  ( .D(n795), .CK(clk), .RN(n25), .Q(\gbuff[20][9] )
         );
  DFFRX1 \gbuff_reg[20][8]  ( .D(n794), .CK(clk), .RN(n24), .Q(\gbuff[20][8] )
         );
  DFFRX1 \gbuff_reg[20][7]  ( .D(n793), .CK(clk), .RN(n17), .Q(\gbuff[20][7] )
         );
  DFFRX1 \gbuff_reg[20][6]  ( .D(n792), .CK(clk), .RN(n18), .Q(\gbuff[20][6] )
         );
  DFFRX1 \gbuff_reg[20][5]  ( .D(n791), .CK(clk), .RN(n25), .Q(\gbuff[20][5] )
         );
  DFFRX1 \gbuff_reg[20][4]  ( .D(n790), .CK(clk), .RN(n19), .Q(\gbuff[20][4] )
         );
  DFFRX1 \gbuff_reg[20][3]  ( .D(n789), .CK(clk), .RN(n24), .Q(\gbuff[20][3] )
         );
  DFFRX1 \gbuff_reg[20][2]  ( .D(n788), .CK(clk), .RN(n17), .Q(\gbuff[20][2] )
         );
  DFFRX1 \gbuff_reg[20][1]  ( .D(n787), .CK(clk), .RN(n20), .Q(\gbuff[20][1] )
         );
  DFFRX1 \gbuff_reg[20][0]  ( .D(n786), .CK(clk), .RN(n23), .Q(\gbuff[20][0] )
         );
  DFFRX1 \gbuff_reg[16][31]  ( .D(n689), .CK(clk), .RN(n19), .Q(
        \gbuff[16][31] ) );
  DFFRX1 \gbuff_reg[16][30]  ( .D(n688), .CK(clk), .RN(n19), .Q(
        \gbuff[16][30] ) );
  DFFRX1 \gbuff_reg[16][29]  ( .D(n687), .CK(clk), .RN(n19), .Q(
        \gbuff[16][29] ) );
  DFFRX1 \gbuff_reg[16][28]  ( .D(n686), .CK(clk), .RN(n26), .Q(
        \gbuff[16][28] ) );
  DFFRX1 \gbuff_reg[16][27]  ( .D(n685), .CK(clk), .RN(n24), .Q(
        \gbuff[16][27] ) );
  DFFRX1 \gbuff_reg[16][26]  ( .D(n684), .CK(clk), .RN(n21), .Q(
        \gbuff[16][26] ) );
  DFFRX1 \gbuff_reg[16][25]  ( .D(n683), .CK(clk), .RN(n24), .Q(
        \gbuff[16][25] ) );
  DFFRX1 \gbuff_reg[16][24]  ( .D(n682), .CK(clk), .RN(n23), .Q(
        \gbuff[16][24] ) );
  DFFRX1 \gbuff_reg[16][23]  ( .D(n681), .CK(clk), .RN(n26), .Q(
        \gbuff[16][23] ) );
  DFFRX1 \gbuff_reg[16][22]  ( .D(n680), .CK(clk), .RN(n20), .Q(
        \gbuff[16][22] ) );
  DFFRX1 \gbuff_reg[16][21]  ( .D(n679), .CK(clk), .RN(n19), .Q(
        \gbuff[16][21] ) );
  DFFRX1 \gbuff_reg[16][20]  ( .D(n678), .CK(clk), .RN(n26), .Q(
        \gbuff[16][20] ) );
  DFFRX1 \gbuff_reg[16][19]  ( .D(n677), .CK(clk), .RN(n21), .Q(
        \gbuff[16][19] ) );
  DFFRX1 \gbuff_reg[16][18]  ( .D(n676), .CK(clk), .RN(n20), .Q(
        \gbuff[16][18] ) );
  DFFRX1 \gbuff_reg[16][17]  ( .D(n675), .CK(clk), .RN(n24), .Q(
        \gbuff[16][17] ) );
  DFFRX1 \gbuff_reg[16][16]  ( .D(n674), .CK(clk), .RN(n17), .Q(
        \gbuff[16][16] ) );
  DFFRX1 \gbuff_reg[16][15]  ( .D(n673), .CK(clk), .RN(n26), .Q(
        \gbuff[16][15] ) );
  DFFRX1 \gbuff_reg[16][14]  ( .D(n672), .CK(clk), .RN(n20), .Q(
        \gbuff[16][14] ) );
  DFFRX1 \gbuff_reg[16][13]  ( .D(n671), .CK(clk), .RN(n26), .Q(
        \gbuff[16][13] ) );
  DFFRX1 \gbuff_reg[16][12]  ( .D(n670), .CK(clk), .RN(n25), .Q(
        \gbuff[16][12] ) );
  DFFRX1 \gbuff_reg[16][11]  ( .D(n669), .CK(clk), .RN(n25), .Q(
        \gbuff[16][11] ) );
  DFFRX1 \gbuff_reg[16][10]  ( .D(n668), .CK(clk), .RN(n21), .Q(
        \gbuff[16][10] ) );
  DFFRX1 \gbuff_reg[16][9]  ( .D(n667), .CK(clk), .RN(n25), .Q(\gbuff[16][9] )
         );
  DFFRX1 \gbuff_reg[16][8]  ( .D(n666), .CK(clk), .RN(n25), .Q(\gbuff[16][8] )
         );
  DFFRX1 \gbuff_reg[16][7]  ( .D(n665), .CK(clk), .RN(n20), .Q(\gbuff[16][7] )
         );
  DFFRX1 \gbuff_reg[16][6]  ( .D(n664), .CK(clk), .RN(n23), .Q(\gbuff[16][6] )
         );
  DFFRX1 \gbuff_reg[16][5]  ( .D(n663), .CK(clk), .RN(n23), .Q(\gbuff[16][5] )
         );
  DFFRX1 \gbuff_reg[16][4]  ( .D(n662), .CK(clk), .RN(n25), .Q(\gbuff[16][4] )
         );
  DFFRX1 \gbuff_reg[16][3]  ( .D(n661), .CK(clk), .RN(n25), .Q(\gbuff[16][3] )
         );
  DFFRX1 \gbuff_reg[16][2]  ( .D(n660), .CK(clk), .RN(n20), .Q(\gbuff[16][2] )
         );
  DFFRX1 \gbuff_reg[16][1]  ( .D(n659), .CK(clk), .RN(n26), .Q(\gbuff[16][1] )
         );
  DFFRX1 \gbuff_reg[16][0]  ( .D(n658), .CK(clk), .RN(n25), .Q(\gbuff[16][0] )
         );
  DFFRX1 \gbuff_reg[12][31]  ( .D(n561), .CK(clk), .RN(n23), .Q(
        \gbuff[12][31] ) );
  DFFRX1 \gbuff_reg[12][30]  ( .D(n560), .CK(clk), .RN(n21), .Q(
        \gbuff[12][30] ) );
  DFFRX1 \gbuff_reg[12][29]  ( .D(n559), .CK(clk), .RN(n23), .Q(
        \gbuff[12][29] ) );
  DFFRX1 \gbuff_reg[12][28]  ( .D(n558), .CK(clk), .RN(n17), .Q(
        \gbuff[12][28] ) );
  DFFRX1 \gbuff_reg[12][27]  ( .D(n557), .CK(clk), .RN(n18), .Q(
        \gbuff[12][27] ) );
  DFFRX1 \gbuff_reg[12][26]  ( .D(n556), .CK(clk), .RN(n17), .Q(
        \gbuff[12][26] ) );
  DFFRX1 \gbuff_reg[12][25]  ( .D(n555), .CK(clk), .RN(n26), .Q(
        \gbuff[12][25] ) );
  DFFRX1 \gbuff_reg[12][24]  ( .D(n554), .CK(clk), .RN(n18), .Q(
        \gbuff[12][24] ) );
  DFFRX1 \gbuff_reg[12][23]  ( .D(n553), .CK(clk), .RN(n23), .Q(
        \gbuff[12][23] ) );
  DFFRX1 \gbuff_reg[12][22]  ( .D(n552), .CK(clk), .RN(n21), .Q(
        \gbuff[12][22] ) );
  DFFRX1 \gbuff_reg[12][21]  ( .D(n551), .CK(clk), .RN(n24), .Q(
        \gbuff[12][21] ) );
  DFFRX1 \gbuff_reg[12][20]  ( .D(n550), .CK(clk), .RN(n23), .Q(
        \gbuff[12][20] ) );
  DFFRX1 \gbuff_reg[12][19]  ( .D(n549), .CK(clk), .RN(n19), .Q(
        \gbuff[12][19] ) );
  DFFRX1 \gbuff_reg[12][18]  ( .D(n548), .CK(clk), .RN(n18), .Q(
        \gbuff[12][18] ) );
  DFFRX1 \gbuff_reg[12][17]  ( .D(n547), .CK(clk), .RN(n21), .Q(
        \gbuff[12][17] ) );
  DFFRX1 \gbuff_reg[12][16]  ( .D(n546), .CK(clk), .RN(n26), .Q(
        \gbuff[12][16] ) );
  DFFRX1 \gbuff_reg[12][15]  ( .D(n545), .CK(clk), .RN(n17), .Q(
        \gbuff[12][15] ) );
  DFFRX1 \gbuff_reg[12][14]  ( .D(n544), .CK(clk), .RN(n25), .Q(
        \gbuff[12][14] ) );
  DFFRX1 \gbuff_reg[12][13]  ( .D(n543), .CK(clk), .RN(n25), .Q(
        \gbuff[12][13] ) );
  DFFRX1 \gbuff_reg[12][12]  ( .D(n542), .CK(clk), .RN(n23), .Q(
        \gbuff[12][12] ) );
  DFFRX1 \gbuff_reg[12][11]  ( .D(n541), .CK(clk), .RN(n19), .Q(
        \gbuff[12][11] ) );
  DFFRX1 \gbuff_reg[12][10]  ( .D(n540), .CK(clk), .RN(n18), .Q(
        \gbuff[12][10] ) );
  DFFRX1 \gbuff_reg[12][9]  ( .D(n539), .CK(clk), .RN(n25), .Q(\gbuff[12][9] )
         );
  DFFRX1 \gbuff_reg[12][8]  ( .D(n538), .CK(clk), .RN(n26), .Q(\gbuff[12][8] )
         );
  DFFRX1 \gbuff_reg[12][7]  ( .D(n537), .CK(clk), .RN(n21), .Q(\gbuff[12][7] )
         );
  DFFRX1 \gbuff_reg[12][6]  ( .D(n536), .CK(clk), .RN(n19), .Q(\gbuff[12][6] )
         );
  DFFRX1 \gbuff_reg[12][5]  ( .D(n535), .CK(clk), .RN(n25), .Q(\gbuff[12][5] )
         );
  DFFRX1 \gbuff_reg[12][4]  ( .D(n534), .CK(clk), .RN(n24), .Q(\gbuff[12][4] )
         );
  DFFRX1 \gbuff_reg[12][3]  ( .D(n533), .CK(clk), .RN(n24), .Q(\gbuff[12][3] )
         );
  DFFRX1 \gbuff_reg[12][2]  ( .D(n532), .CK(clk), .RN(n21), .Q(\gbuff[12][2] )
         );
  DFFRX1 \gbuff_reg[12][1]  ( .D(n531), .CK(clk), .RN(n17), .Q(\gbuff[12][1] )
         );
  DFFRX1 \gbuff_reg[12][0]  ( .D(n530), .CK(clk), .RN(n20), .Q(\gbuff[12][0] )
         );
  DFFRX1 \gbuff_reg[8][31]  ( .D(n433), .CK(clk), .RN(n21), .Q(\gbuff[8][31] )
         );
  DFFRX1 \gbuff_reg[8][30]  ( .D(n432), .CK(clk), .RN(n19), .Q(\gbuff[8][30] )
         );
  DFFRX1 \gbuff_reg[8][29]  ( .D(n431), .CK(clk), .RN(n17), .Q(\gbuff[8][29] )
         );
  DFFRX1 \gbuff_reg[8][28]  ( .D(n430), .CK(clk), .RN(n26), .Q(\gbuff[8][28] )
         );
  DFFRX1 \gbuff_reg[8][27]  ( .D(n429), .CK(clk), .RN(n20), .Q(\gbuff[8][27] )
         );
  DFFRX1 \gbuff_reg[8][26]  ( .D(n428), .CK(clk), .RN(n19), .Q(\gbuff[8][26] )
         );
  DFFRX1 \gbuff_reg[8][25]  ( .D(n427), .CK(clk), .RN(n26), .Q(\gbuff[8][25] )
         );
  DFFRX1 \gbuff_reg[8][24]  ( .D(n426), .CK(clk), .RN(n24), .Q(\gbuff[8][24] )
         );
  DFFRX1 \gbuff_reg[8][23]  ( .D(n425), .CK(clk), .RN(n26), .Q(\gbuff[8][23] )
         );
  DFFRX1 \gbuff_reg[8][22]  ( .D(n424), .CK(clk), .RN(n26), .Q(\gbuff[8][22] )
         );
  DFFRX1 \gbuff_reg[8][21]  ( .D(n423), .CK(clk), .RN(n26), .Q(\gbuff[8][21] )
         );
  DFFRX1 \gbuff_reg[8][20]  ( .D(n422), .CK(clk), .RN(n19), .Q(\gbuff[8][20] )
         );
  DFFRX1 \gbuff_reg[8][19]  ( .D(n421), .CK(clk), .RN(n20), .Q(\gbuff[8][19] )
         );
  DFFRX1 \gbuff_reg[8][18]  ( .D(n420), .CK(clk), .RN(n17), .Q(\gbuff[8][18] )
         );
  DFFRX1 \gbuff_reg[8][17]  ( .D(n419), .CK(clk), .RN(n23), .Q(\gbuff[8][17] )
         );
  DFFRX1 \gbuff_reg[8][16]  ( .D(n418), .CK(clk), .RN(n24), .Q(\gbuff[8][16] )
         );
  DFFRX1 \gbuff_reg[8][15]  ( .D(n417), .CK(clk), .RN(n18), .Q(\gbuff[8][15] )
         );
  DFFRX1 \gbuff_reg[8][14]  ( .D(n416), .CK(clk), .RN(n23), .Q(\gbuff[8][14] )
         );
  DFFRX1 \gbuff_reg[8][13]  ( .D(n415), .CK(clk), .RN(n26), .Q(\gbuff[8][13] )
         );
  DFFRX1 \gbuff_reg[8][12]  ( .D(n414), .CK(clk), .RN(n18), .Q(\gbuff[8][12] )
         );
  DFFRX1 \gbuff_reg[8][11]  ( .D(n413), .CK(clk), .RN(n25), .Q(\gbuff[8][11] )
         );
  DFFRX1 \gbuff_reg[8][10]  ( .D(n412), .CK(clk), .RN(n18), .Q(\gbuff[8][10] )
         );
  DFFRX1 \gbuff_reg[8][9]  ( .D(n411), .CK(clk), .RN(n24), .Q(\gbuff[8][9] )
         );
  DFFRX1 \gbuff_reg[8][8]  ( .D(n410), .CK(clk), .RN(n21), .Q(\gbuff[8][8] )
         );
  DFFRX1 \gbuff_reg[8][7]  ( .D(n409), .CK(clk), .RN(n18), .Q(\gbuff[8][7] )
         );
  DFFRX1 \gbuff_reg[8][6]  ( .D(n408), .CK(clk), .RN(n23), .Q(\gbuff[8][6] )
         );
  DFFRX1 \gbuff_reg[8][5]  ( .D(n407), .CK(clk), .RN(n18), .Q(\gbuff[8][5] )
         );
  DFFRX1 \gbuff_reg[8][4]  ( .D(n406), .CK(clk), .RN(n25), .Q(\gbuff[8][4] )
         );
  DFFRX1 \gbuff_reg[8][3]  ( .D(n405), .CK(clk), .RN(n17), .Q(\gbuff[8][3] )
         );
  DFFRX1 \gbuff_reg[8][2]  ( .D(n404), .CK(clk), .RN(n20), .Q(\gbuff[8][2] )
         );
  DFFRX1 \gbuff_reg[8][1]  ( .D(n403), .CK(clk), .RN(n19), .Q(\gbuff[8][1] )
         );
  DFFRX1 \gbuff_reg[8][0]  ( .D(n402), .CK(clk), .RN(n17), .Q(\gbuff[8][0] )
         );
  DFFRX1 \gbuff_reg[4][31]  ( .D(n305), .CK(clk), .RN(n23), .Q(\gbuff[4][31] )
         );
  DFFRX1 \gbuff_reg[4][30]  ( .D(n304), .CK(clk), .RN(n24), .Q(\gbuff[4][30] )
         );
  DFFRX1 \gbuff_reg[4][29]  ( .D(n303), .CK(clk), .RN(n24), .Q(\gbuff[4][29] )
         );
  DFFRX1 \gbuff_reg[4][28]  ( .D(n302), .CK(clk), .RN(n21), .Q(\gbuff[4][28] )
         );
  DFFRX1 \gbuff_reg[4][27]  ( .D(n301), .CK(clk), .RN(n17), .Q(\gbuff[4][27] )
         );
  DFFRX1 \gbuff_reg[4][26]  ( .D(n300), .CK(clk), .RN(n24), .Q(\gbuff[4][26] )
         );
  DFFRX1 \gbuff_reg[4][25]  ( .D(n299), .CK(clk), .RN(n19), .Q(\gbuff[4][25] )
         );
  DFFRX1 \gbuff_reg[4][24]  ( .D(n298), .CK(clk), .RN(n17), .Q(\gbuff[4][24] )
         );
  DFFRX1 \gbuff_reg[4][23]  ( .D(n297), .CK(clk), .RN(n24), .Q(\gbuff[4][23] )
         );
  DFFRX1 \gbuff_reg[4][22]  ( .D(n296), .CK(clk), .RN(n25), .Q(\gbuff[4][22] )
         );
  DFFRX1 \gbuff_reg[4][21]  ( .D(n295), .CK(clk), .RN(n24), .Q(\gbuff[4][21] )
         );
  DFFRX1 \gbuff_reg[4][20]  ( .D(n294), .CK(clk), .RN(n17), .Q(\gbuff[4][20] )
         );
  DFFRX1 \gbuff_reg[4][19]  ( .D(n293), .CK(clk), .RN(n19), .Q(\gbuff[4][19] )
         );
  DFFRX1 \gbuff_reg[4][18]  ( .D(n292), .CK(clk), .RN(n19), .Q(\gbuff[4][18] )
         );
  DFFRX1 \gbuff_reg[4][17]  ( .D(n291), .CK(clk), .RN(n18), .Q(\gbuff[4][17] )
         );
  DFFRX1 \gbuff_reg[4][16]  ( .D(n290), .CK(clk), .RN(n19), .Q(\gbuff[4][16] )
         );
  DFFRX1 \gbuff_reg[4][15]  ( .D(n289), .CK(clk), .RN(n24), .Q(\gbuff[4][15] )
         );
  DFFRX1 \gbuff_reg[4][14]  ( .D(n288), .CK(clk), .RN(n25), .Q(\gbuff[4][14] )
         );
  DFFRX1 \gbuff_reg[4][13]  ( .D(n287), .CK(clk), .RN(n20), .Q(\gbuff[4][13] )
         );
  DFFRX1 \gbuff_reg[4][12]  ( .D(n286), .CK(clk), .RN(n24), .Q(\gbuff[4][12] )
         );
  DFFRX1 \gbuff_reg[4][11]  ( .D(n285), .CK(clk), .RN(n26), .Q(\gbuff[4][11] )
         );
  DFFRX1 \gbuff_reg[4][10]  ( .D(n284), .CK(clk), .RN(n23), .Q(\gbuff[4][10] )
         );
  DFFRX1 \gbuff_reg[4][9]  ( .D(n283), .CK(clk), .RN(n24), .Q(\gbuff[4][9] )
         );
  DFFRX1 \gbuff_reg[4][8]  ( .D(n282), .CK(clk), .RN(n18), .Q(\gbuff[4][8] )
         );
  DFFRX1 \gbuff_reg[4][7]  ( .D(n281), .CK(clk), .RN(n21), .Q(\gbuff[4][7] )
         );
  DFFRX1 \gbuff_reg[4][6]  ( .D(n280), .CK(clk), .RN(n17), .Q(\gbuff[4][6] )
         );
  DFFRX1 \gbuff_reg[4][5]  ( .D(n279), .CK(clk), .RN(n17), .Q(\gbuff[4][5] )
         );
  DFFRX1 \gbuff_reg[4][4]  ( .D(n278), .CK(clk), .RN(n20), .Q(\gbuff[4][4] )
         );
  DFFRX1 \gbuff_reg[4][3]  ( .D(n277), .CK(clk), .RN(n26), .Q(\gbuff[4][3] )
         );
  DFFRX1 \gbuff_reg[4][2]  ( .D(n276), .CK(clk), .RN(n26), .Q(\gbuff[4][2] )
         );
  DFFRX1 \gbuff_reg[4][1]  ( .D(n275), .CK(clk), .RN(n21), .Q(\gbuff[4][1] )
         );
  DFFRX1 \gbuff_reg[4][0]  ( .D(n274), .CK(clk), .RN(n18), .Q(\gbuff[4][0] )
         );
  DFFRX1 \gbuff_reg[0][31]  ( .D(n177), .CK(clk), .RN(n25), .Q(\gbuff[0][31] )
         );
  DFFRX1 \gbuff_reg[0][30]  ( .D(n176), .CK(clk), .RN(n26), .Q(\gbuff[0][30] )
         );
  DFFRX1 \gbuff_reg[0][29]  ( .D(n175), .CK(clk), .RN(n17), .Q(\gbuff[0][29] )
         );
  DFFRX1 \gbuff_reg[0][28]  ( .D(n174), .CK(clk), .RN(n20), .Q(\gbuff[0][28] )
         );
  DFFRX1 \gbuff_reg[0][27]  ( .D(n173), .CK(clk), .RN(n20), .Q(\gbuff[0][27] )
         );
  DFFRX1 \gbuff_reg[0][26]  ( .D(n172), .CK(clk), .RN(n20), .Q(\gbuff[0][26] )
         );
  DFFRX1 \gbuff_reg[0][25]  ( .D(n171), .CK(clk), .RN(n17), .Q(\gbuff[0][25] )
         );
  DFFRX1 \gbuff_reg[0][24]  ( .D(n170), .CK(clk), .RN(n23), .Q(\gbuff[0][24] )
         );
  DFFRX1 \gbuff_reg[0][23]  ( .D(n169), .CK(clk), .RN(n25), .Q(\gbuff[0][23] )
         );
  DFFRX1 \gbuff_reg[0][22]  ( .D(n168), .CK(clk), .RN(n26), .Q(\gbuff[0][22] )
         );
  DFFRX1 \gbuff_reg[0][21]  ( .D(n167), .CK(clk), .RN(n21), .Q(\gbuff[0][21] )
         );
  DFFRX1 \gbuff_reg[0][20]  ( .D(n166), .CK(clk), .RN(n26), .Q(\gbuff[0][20] )
         );
  DFFRX1 \gbuff_reg[0][19]  ( .D(n165), .CK(clk), .RN(n23), .Q(\gbuff[0][19] )
         );
  DFFRX1 \gbuff_reg[0][18]  ( .D(n164), .CK(clk), .RN(n21), .Q(\gbuff[0][18] )
         );
  DFFRX1 \gbuff_reg[0][17]  ( .D(n163), .CK(clk), .RN(n23), .Q(\gbuff[0][17] )
         );
  DFFRX1 \gbuff_reg[0][16]  ( .D(n162), .CK(clk), .RN(n20), .Q(\gbuff[0][16] )
         );
  DFFRX1 \gbuff_reg[0][15]  ( .D(n161), .CK(clk), .RN(n18), .Q(\gbuff[0][15] )
         );
  DFFRX1 \gbuff_reg[0][14]  ( .D(n160), .CK(clk), .RN(n18), .Q(\gbuff[0][14] )
         );
  DFFRX1 \gbuff_reg[0][13]  ( .D(n159), .CK(clk), .RN(n18), .Q(\gbuff[0][13] )
         );
  DFFRX1 \gbuff_reg[0][12]  ( .D(n158), .CK(clk), .RN(n18), .Q(\gbuff[0][12] )
         );
  DFFRX1 \gbuff_reg[0][11]  ( .D(n157), .CK(clk), .RN(n23), .Q(\gbuff[0][11] )
         );
  DFFRX1 \gbuff_reg[0][10]  ( .D(n156), .CK(clk), .RN(n25), .Q(\gbuff[0][10] )
         );
  DFFRX1 \gbuff_reg[0][9]  ( .D(n155), .CK(clk), .RN(n20), .Q(\gbuff[0][9] )
         );
  DFFRX1 \gbuff_reg[0][8]  ( .D(n154), .CK(clk), .RN(n20), .Q(\gbuff[0][8] )
         );
  DFFRX1 \gbuff_reg[0][7]  ( .D(n153), .CK(clk), .RN(n19), .Q(\gbuff[0][7] )
         );
  DFFRX1 \gbuff_reg[0][6]  ( .D(n152), .CK(clk), .RN(n24), .Q(\gbuff[0][6] )
         );
  DFFRX1 \gbuff_reg[0][5]  ( .D(n151), .CK(clk), .RN(n18), .Q(\gbuff[0][5] )
         );
  DFFRX1 \gbuff_reg[0][4]  ( .D(n150), .CK(clk), .RN(n18), .Q(\gbuff[0][4] )
         );
  DFFRX1 \gbuff_reg[0][3]  ( .D(n149), .CK(clk), .RN(n17), .Q(\gbuff[0][3] )
         );
  DFFRX1 \gbuff_reg[0][2]  ( .D(n148), .CK(clk), .RN(n23), .Q(\gbuff[0][2] )
         );
  DFFRX1 \gbuff_reg[0][1]  ( .D(n147), .CK(clk), .RN(n20), .Q(\gbuff[0][1] )
         );
  DFFRX1 \gbuff_reg[0][0]  ( .D(n146), .CK(clk), .RN(n25), .Q(\gbuff[0][0] )
         );
  DFFRX1 \gbuff_reg[31][31]  ( .D(n1169), .CK(clk), .RN(n19), .Q(
        \gbuff[31][31] ) );
  DFFRX1 \gbuff_reg[31][30]  ( .D(n1168), .CK(clk), .RN(n24), .Q(
        \gbuff[31][30] ) );
  DFFRX1 \gbuff_reg[31][29]  ( .D(n1167), .CK(clk), .RN(n19), .Q(
        \gbuff[31][29] ) );
  DFFRX1 \gbuff_reg[31][28]  ( .D(n1166), .CK(clk), .RN(n17), .Q(
        \gbuff[31][28] ) );
  DFFRX1 \gbuff_reg[31][27]  ( .D(n1165), .CK(clk), .RN(n21), .Q(
        \gbuff[31][27] ) );
  DFFRX1 \gbuff_reg[31][26]  ( .D(n1164), .CK(clk), .RN(n25), .Q(
        \gbuff[31][26] ) );
  DFFRX1 \gbuff_reg[31][25]  ( .D(n1163), .CK(clk), .RN(n17), .Q(
        \gbuff[31][25] ) );
  DFFRX1 \gbuff_reg[31][24]  ( .D(n1162), .CK(clk), .RN(n21), .Q(
        \gbuff[31][24] ) );
  DFFRX1 \gbuff_reg[31][23]  ( .D(n1161), .CK(clk), .RN(n24), .Q(
        \gbuff[31][23] ) );
  DFFRX1 \gbuff_reg[31][22]  ( .D(n1160), .CK(clk), .RN(n20), .Q(
        \gbuff[31][22] ) );
  DFFRX1 \gbuff_reg[31][21]  ( .D(n1159), .CK(clk), .RN(n20), .Q(
        \gbuff[31][21] ) );
  DFFRX1 \gbuff_reg[31][20]  ( .D(n1158), .CK(clk), .RN(n17), .Q(
        \gbuff[31][20] ) );
  DFFRX1 \gbuff_reg[31][19]  ( .D(n1157), .CK(clk), .RN(n21), .Q(
        \gbuff[31][19] ) );
  DFFRX1 \gbuff_reg[31][18]  ( .D(n1156), .CK(clk), .RN(n23), .Q(
        \gbuff[31][18] ) );
  DFFRX1 \gbuff_reg[31][17]  ( .D(n1155), .CK(clk), .RN(n18), .Q(
        \gbuff[31][17] ) );
  DFFRX1 \gbuff_reg[31][16]  ( .D(n1154), .CK(clk), .RN(n21), .Q(
        \gbuff[31][16] ) );
  DFFRX1 \gbuff_reg[31][15]  ( .D(n1153), .CK(clk), .RN(n20), .Q(
        \gbuff[31][15] ) );
  DFFRX1 \gbuff_reg[31][14]  ( .D(n1152), .CK(clk), .RN(n17), .Q(
        \gbuff[31][14] ) );
  DFFRX1 \gbuff_reg[31][13]  ( .D(n1151), .CK(clk), .RN(n20), .Q(
        \gbuff[31][13] ) );
  DFFRX1 \gbuff_reg[31][12]  ( .D(n1150), .CK(clk), .RN(n21), .Q(
        \gbuff[31][12] ) );
  DFFRX1 \gbuff_reg[31][11]  ( .D(n1149), .CK(clk), .RN(n26), .Q(
        \gbuff[31][11] ) );
  DFFRX1 \gbuff_reg[31][10]  ( .D(n1148), .CK(clk), .RN(n21), .Q(
        \gbuff[31][10] ) );
  DFFRX1 \gbuff_reg[31][9]  ( .D(n1147), .CK(clk), .RN(n18), .Q(\gbuff[31][9] ) );
  DFFRX1 \gbuff_reg[31][8]  ( .D(n1146), .CK(clk), .RN(n26), .Q(\gbuff[31][8] ) );
  DFFRX1 \gbuff_reg[31][7]  ( .D(n1145), .CK(clk), .RN(n20), .Q(\gbuff[31][7] ) );
  DFFRX1 \gbuff_reg[31][6]  ( .D(n1144), .CK(clk), .RN(n17), .Q(\gbuff[31][6] ) );
  DFFRX1 \gbuff_reg[31][5]  ( .D(n1143), .CK(clk), .RN(n23), .Q(\gbuff[31][5] ) );
  DFFRX1 \gbuff_reg[31][4]  ( .D(n1142), .CK(clk), .RN(n24), .Q(\gbuff[31][4] ) );
  DFFRX1 \gbuff_reg[31][3]  ( .D(n1141), .CK(clk), .RN(n18), .Q(\gbuff[31][3] ) );
  DFFRX1 \gbuff_reg[31][2]  ( .D(n1140), .CK(clk), .RN(n19), .Q(\gbuff[31][2] ) );
  DFFRX1 \gbuff_reg[31][1]  ( .D(n1139), .CK(clk), .RN(n25), .Q(\gbuff[31][1] ) );
  DFFRX1 \gbuff_reg[31][0]  ( .D(n1138), .CK(clk), .RN(n19), .Q(\gbuff[31][0] ) );
  DFFRX1 \gbuff_reg[27][31]  ( .D(n1041), .CK(clk), .RN(n25), .Q(
        \gbuff[27][31] ) );
  DFFRX1 \gbuff_reg[27][30]  ( .D(n1040), .CK(clk), .RN(n21), .Q(
        \gbuff[27][30] ) );
  DFFRX1 \gbuff_reg[27][29]  ( .D(n1039), .CK(clk), .RN(n21), .Q(
        \gbuff[27][29] ) );
  DFFRX1 \gbuff_reg[27][28]  ( .D(n1038), .CK(clk), .RN(n24), .Q(
        \gbuff[27][28] ) );
  DFFRX1 \gbuff_reg[27][27]  ( .D(n1037), .CK(clk), .RN(n18), .Q(
        \gbuff[27][27] ) );
  DFFRX1 \gbuff_reg[27][26]  ( .D(n1036), .CK(clk), .RN(n19), .Q(
        \gbuff[27][26] ) );
  DFFRX1 \gbuff_reg[27][25]  ( .D(n1035), .CK(clk), .RN(n17), .Q(
        \gbuff[27][25] ) );
  DFFRX1 \gbuff_reg[27][24]  ( .D(n1034), .CK(clk), .RN(n19), .Q(
        \gbuff[27][24] ) );
  DFFRX1 \gbuff_reg[27][23]  ( .D(n1033), .CK(clk), .RN(n17), .Q(
        \gbuff[27][23] ) );
  DFFRX1 \gbuff_reg[27][22]  ( .D(n1032), .CK(clk), .RN(n18), .Q(
        \gbuff[27][22] ) );
  DFFRX1 \gbuff_reg[27][21]  ( .D(n1031), .CK(clk), .RN(n21), .Q(
        \gbuff[27][21] ) );
  DFFRX1 \gbuff_reg[27][20]  ( .D(n1030), .CK(clk), .RN(n20), .Q(
        \gbuff[27][20] ) );
  DFFRX1 \gbuff_reg[27][19]  ( .D(n1029), .CK(clk), .RN(n23), .Q(
        \gbuff[27][19] ) );
  DFFRX1 \gbuff_reg[27][18]  ( .D(n1028), .CK(clk), .RN(n25), .Q(
        \gbuff[27][18] ) );
  DFFRX1 \gbuff_reg[27][17]  ( .D(n1027), .CK(clk), .RN(n21), .Q(
        \gbuff[27][17] ) );
  DFFRX1 \gbuff_reg[27][16]  ( .D(n1026), .CK(clk), .RN(n24), .Q(
        \gbuff[27][16] ) );
  DFFRX1 \gbuff_reg[27][15]  ( .D(n1025), .CK(clk), .RN(n17), .Q(
        \gbuff[27][15] ) );
  DFFRX1 \gbuff_reg[27][14]  ( .D(n1024), .CK(clk), .RN(n18), .Q(
        \gbuff[27][14] ) );
  DFFRX1 \gbuff_reg[27][13]  ( .D(n1023), .CK(clk), .RN(n25), .Q(
        \gbuff[27][13] ) );
  DFFRX1 \gbuff_reg[27][12]  ( .D(n1022), .CK(clk), .RN(n18), .Q(
        \gbuff[27][12] ) );
  DFFRX1 \gbuff_reg[27][11]  ( .D(n1021), .CK(clk), .RN(n24), .Q(
        \gbuff[27][11] ) );
  DFFRX1 \gbuff_reg[27][10]  ( .D(n1020), .CK(clk), .RN(n26), .Q(
        \gbuff[27][10] ) );
  DFFRX1 \gbuff_reg[27][9]  ( .D(n1019), .CK(clk), .RN(n18), .Q(\gbuff[27][9] ) );
  DFFRX1 \gbuff_reg[27][8]  ( .D(n1018), .CK(clk), .RN(n23), .Q(\gbuff[27][8] ) );
  DFFRX1 \gbuff_reg[27][7]  ( .D(n1017), .CK(clk), .RN(n19), .Q(\gbuff[27][7] ) );
  DFFRX1 \gbuff_reg[27][6]  ( .D(n1016), .CK(clk), .RN(n19), .Q(\gbuff[27][6] ) );
  DFFRX1 \gbuff_reg[27][5]  ( .D(n1015), .CK(clk), .RN(n19), .Q(\gbuff[27][5] ) );
  DFFRX1 \gbuff_reg[27][4]  ( .D(n1014), .CK(clk), .RN(n26), .Q(\gbuff[27][4] ) );
  DFFRX1 \gbuff_reg[27][3]  ( .D(n1013), .CK(clk), .RN(n24), .Q(\gbuff[27][3] ) );
  DFFRX1 \gbuff_reg[27][2]  ( .D(n1012), .CK(clk), .RN(n21), .Q(\gbuff[27][2] ) );
  DFFRX1 \gbuff_reg[27][1]  ( .D(n1011), .CK(clk), .RN(n24), .Q(\gbuff[27][1] ) );
  DFFRX1 \gbuff_reg[27][0]  ( .D(n1010), .CK(clk), .RN(n23), .Q(\gbuff[27][0] ) );
  DFFRX1 \gbuff_reg[23][31]  ( .D(n913), .CK(clk), .RN(n26), .Q(
        \gbuff[23][31] ) );
  DFFRX1 \gbuff_reg[23][30]  ( .D(n912), .CK(clk), .RN(n20), .Q(
        \gbuff[23][30] ) );
  DFFRX1 \gbuff_reg[23][29]  ( .D(n911), .CK(clk), .RN(n19), .Q(
        \gbuff[23][29] ) );
  DFFRX1 \gbuff_reg[23][28]  ( .D(n910), .CK(clk), .RN(n19), .Q(
        \gbuff[23][28] ) );
  DFFRX1 \gbuff_reg[23][27]  ( .D(n909), .CK(clk), .RN(n21), .Q(
        \gbuff[23][27] ) );
  DFFRX1 \gbuff_reg[23][26]  ( .D(n908), .CK(clk), .RN(n19), .Q(
        \gbuff[23][26] ) );
  DFFRX1 \gbuff_reg[23][25]  ( .D(n907), .CK(clk), .RN(n20), .Q(
        \gbuff[23][25] ) );
  DFFRX1 \gbuff_reg[23][24]  ( .D(n906), .CK(clk), .RN(n17), .Q(
        \gbuff[23][24] ) );
  DFFRX1 \gbuff_reg[23][23]  ( .D(n905), .CK(clk), .RN(n26), .Q(
        \gbuff[23][23] ) );
  DFFRX1 \gbuff_reg[23][22]  ( .D(n904), .CK(clk), .RN(n20), .Q(
        \gbuff[23][22] ) );
  DFFRX1 \gbuff_reg[23][21]  ( .D(n903), .CK(clk), .RN(n26), .Q(
        \gbuff[23][21] ) );
  DFFRX1 \gbuff_reg[23][20]  ( .D(n902), .CK(clk), .RN(n17), .Q(
        \gbuff[23][20] ) );
  DFFRX1 \gbuff_reg[23][19]  ( .D(n901), .CK(clk), .RN(n25), .Q(
        \gbuff[23][19] ) );
  DFFRX1 \gbuff_reg[23][18]  ( .D(n900), .CK(clk), .RN(n23), .Q(
        \gbuff[23][18] ) );
  DFFRX1 \gbuff_reg[23][17]  ( .D(n899), .CK(clk), .RN(n26), .Q(
        \gbuff[23][17] ) );
  DFFRX1 \gbuff_reg[23][16]  ( .D(n898), .CK(clk), .RN(n25), .Q(
        \gbuff[23][16] ) );
  DFFRX1 \gbuff_reg[23][15]  ( .D(n897), .CK(clk), .RN(n20), .Q(
        \gbuff[23][15] ) );
  DFFRX1 \gbuff_reg[23][14]  ( .D(n896), .CK(clk), .RN(n23), .Q(
        \gbuff[23][14] ) );
  DFFRX1 \gbuff_reg[23][13]  ( .D(n895), .CK(clk), .RN(n23), .Q(
        \gbuff[23][13] ) );
  DFFRX1 \gbuff_reg[23][12]  ( .D(n894), .CK(clk), .RN(n25), .Q(
        \gbuff[23][12] ) );
  DFFRX1 \gbuff_reg[23][11]  ( .D(n893), .CK(clk), .RN(n25), .Q(
        \gbuff[23][11] ) );
  DFFRX1 \gbuff_reg[23][10]  ( .D(n892), .CK(clk), .RN(n20), .Q(
        \gbuff[23][10] ) );
  DFFRX1 \gbuff_reg[23][9]  ( .D(n891), .CK(clk), .RN(n26), .Q(\gbuff[23][9] )
         );
  DFFRX1 \gbuff_reg[23][8]  ( .D(n890), .CK(clk), .RN(n25), .Q(\gbuff[23][8] )
         );
  DFFRX1 \gbuff_reg[23][7]  ( .D(n889), .CK(clk), .RN(n23), .Q(\gbuff[23][7] )
         );
  DFFRX1 \gbuff_reg[23][6]  ( .D(n888), .CK(clk), .RN(n21), .Q(\gbuff[23][6] )
         );
  DFFRX1 \gbuff_reg[23][5]  ( .D(n887), .CK(clk), .RN(n23), .Q(\gbuff[23][5] )
         );
  DFFRX1 \gbuff_reg[23][4]  ( .D(n886), .CK(clk), .RN(n21), .Q(\gbuff[23][4] )
         );
  DFFRX1 \gbuff_reg[23][3]  ( .D(n885), .CK(clk), .RN(n18), .Q(\gbuff[23][3] )
         );
  DFFRX1 \gbuff_reg[23][2]  ( .D(n884), .CK(clk), .RN(n26), .Q(\gbuff[23][2] )
         );
  DFFRX1 \gbuff_reg[23][1]  ( .D(n883), .CK(clk), .RN(n19), .Q(\gbuff[23][1] )
         );
  DFFRX1 \gbuff_reg[23][0]  ( .D(n882), .CK(clk), .RN(n18), .Q(\gbuff[23][0] )
         );
  DFFRX1 \gbuff_reg[19][31]  ( .D(n785), .CK(clk), .RN(n23), .Q(
        \gbuff[19][31] ) );
  DFFRX1 \gbuff_reg[19][30]  ( .D(n784), .CK(clk), .RN(n21), .Q(
        \gbuff[19][30] ) );
  DFFRX1 \gbuff_reg[19][29]  ( .D(n783), .CK(clk), .RN(n24), .Q(
        \gbuff[19][29] ) );
  DFFRX1 \gbuff_reg[19][28]  ( .D(n782), .CK(clk), .RN(n20), .Q(
        \gbuff[19][28] ) );
  DFFRX1 \gbuff_reg[19][27]  ( .D(n781), .CK(clk), .RN(n19), .Q(
        \gbuff[19][27] ) );
  DFFRX1 \gbuff_reg[19][26]  ( .D(n780), .CK(clk), .RN(n24), .Q(
        \gbuff[19][26] ) );
  DFFRX1 \gbuff_reg[19][25]  ( .D(n779), .CK(clk), .RN(n20), .Q(
        \gbuff[19][25] ) );
  DFFRX1 \gbuff_reg[19][24]  ( .D(n778), .CK(clk), .RN(n26), .Q(
        \gbuff[19][24] ) );
  DFFRX1 \gbuff_reg[19][23]  ( .D(n777), .CK(clk), .RN(n17), .Q(
        \gbuff[19][23] ) );
  DFFRX1 \gbuff_reg[19][22]  ( .D(n776), .CK(clk), .RN(n25), .Q(
        \gbuff[19][22] ) );
  DFFRX1 \gbuff_reg[19][21]  ( .D(n775), .CK(clk), .RN(n25), .Q(
        \gbuff[19][21] ) );
  DFFRX1 \gbuff_reg[19][20]  ( .D(n774), .CK(clk), .RN(n23), .Q(
        \gbuff[19][20] ) );
  DFFRX1 \gbuff_reg[19][19]  ( .D(n773), .CK(clk), .RN(n19), .Q(
        \gbuff[19][19] ) );
  DFFRX1 \gbuff_reg[19][18]  ( .D(n772), .CK(clk), .RN(n18), .Q(
        \gbuff[19][18] ) );
  DFFRX1 \gbuff_reg[19][17]  ( .D(n771), .CK(clk), .RN(n25), .Q(
        \gbuff[19][17] ) );
  DFFRX1 \gbuff_reg[19][16]  ( .D(n770), .CK(clk), .RN(n26), .Q(
        \gbuff[19][16] ) );
  DFFRX1 \gbuff_reg[19][15]  ( .D(n769), .CK(clk), .RN(n21), .Q(
        \gbuff[19][15] ) );
  DFFRX1 \gbuff_reg[19][14]  ( .D(n768), .CK(clk), .RN(n19), .Q(
        \gbuff[19][14] ) );
  DFFRX1 \gbuff_reg[19][13]  ( .D(n767), .CK(clk), .RN(n25), .Q(
        \gbuff[19][13] ) );
  DFFRX1 \gbuff_reg[19][12]  ( .D(n766), .CK(clk), .RN(n23), .Q(
        \gbuff[19][12] ) );
  DFFRX1 \gbuff_reg[19][11]  ( .D(n765), .CK(clk), .RN(n24), .Q(
        \gbuff[19][11] ) );
  DFFRX1 \gbuff_reg[19][10]  ( .D(n764), .CK(clk), .RN(n23), .Q(
        \gbuff[19][10] ) );
  DFFRX1 \gbuff_reg[19][9]  ( .D(n763), .CK(clk), .RN(n21), .Q(\gbuff[19][9] )
         );
  DFFRX1 \gbuff_reg[19][8]  ( .D(n762), .CK(clk), .RN(n20), .Q(\gbuff[19][8] )
         );
  DFFRX1 \gbuff_reg[19][7]  ( .D(n761), .CK(clk), .RN(n21), .Q(\gbuff[19][7] )
         );
  DFFRX1 \gbuff_reg[19][6]  ( .D(n760), .CK(clk), .RN(n19), .Q(\gbuff[19][6] )
         );
  DFFRX1 \gbuff_reg[19][5]  ( .D(n759), .CK(clk), .RN(n17), .Q(\gbuff[19][5] )
         );
  DFFRX1 \gbuff_reg[19][4]  ( .D(n758), .CK(clk), .RN(n18), .Q(\gbuff[19][4] )
         );
  DFFRX1 \gbuff_reg[19][3]  ( .D(n757), .CK(clk), .RN(n20), .Q(\gbuff[19][3] )
         );
  DFFRX1 \gbuff_reg[19][2]  ( .D(n756), .CK(clk), .RN(n25), .Q(\gbuff[19][2] )
         );
  DFFRX1 \gbuff_reg[19][1]  ( .D(n755), .CK(clk), .RN(n24), .Q(\gbuff[19][1] )
         );
  DFFRX1 \gbuff_reg[19][0]  ( .D(n754), .CK(clk), .RN(n24), .Q(\gbuff[19][0] )
         );
  DFFRX1 \gbuff_reg[15][31]  ( .D(n657), .CK(clk), .RN(n26), .Q(
        \gbuff[15][31] ) );
  DFFRX1 \gbuff_reg[15][30]  ( .D(n656), .CK(clk), .RN(n26), .Q(
        \gbuff[15][30] ) );
  DFFRX1 \gbuff_reg[15][29]  ( .D(n655), .CK(clk), .RN(n26), .Q(
        \gbuff[15][29] ) );
  DFFRX1 \gbuff_reg[15][28]  ( .D(n654), .CK(clk), .RN(n19), .Q(
        \gbuff[15][28] ) );
  DFFRX1 \gbuff_reg[15][27]  ( .D(n653), .CK(clk), .RN(n20), .Q(
        \gbuff[15][27] ) );
  DFFRX1 \gbuff_reg[15][26]  ( .D(n652), .CK(clk), .RN(n17), .Q(
        \gbuff[15][26] ) );
  DFFRX1 \gbuff_reg[15][25]  ( .D(n651), .CK(clk), .RN(n23), .Q(
        \gbuff[15][25] ) );
  DFFRX1 \gbuff_reg[15][24]  ( .D(n650), .CK(clk), .RN(n24), .Q(
        \gbuff[15][24] ) );
  DFFRX1 \gbuff_reg[15][23]  ( .D(n649), .CK(clk), .RN(n18), .Q(
        \gbuff[15][23] ) );
  DFFRX1 \gbuff_reg[15][22]  ( .D(n648), .CK(clk), .RN(n23), .Q(
        \gbuff[15][22] ) );
  DFFRX1 \gbuff_reg[15][21]  ( .D(n647), .CK(clk), .RN(n26), .Q(
        \gbuff[15][21] ) );
  DFFRX1 \gbuff_reg[15][20]  ( .D(n646), .CK(clk), .RN(n19), .Q(
        \gbuff[15][20] ) );
  DFFRX1 \gbuff_reg[15][19]  ( .D(n645), .CK(clk), .RN(n25), .Q(
        \gbuff[15][19] ) );
  DFFRX1 \gbuff_reg[15][18]  ( .D(n644), .CK(clk), .RN(n24), .Q(
        \gbuff[15][18] ) );
  DFFRX1 \gbuff_reg[15][17]  ( .D(n643), .CK(clk), .RN(n23), .Q(
        \gbuff[15][17] ) );
  DFFRX1 \gbuff_reg[15][16]  ( .D(n642), .CK(clk), .RN(n21), .Q(
        \gbuff[15][16] ) );
  DFFRX1 \gbuff_reg[15][15]  ( .D(n641), .CK(clk), .RN(n18), .Q(
        \gbuff[15][15] ) );
  DFFRX1 \gbuff_reg[15][14]  ( .D(n640), .CK(clk), .RN(n23), .Q(
        \gbuff[15][14] ) );
  DFFRX1 \gbuff_reg[15][13]  ( .D(n639), .CK(clk), .RN(n18), .Q(
        \gbuff[15][13] ) );
  DFFRX1 \gbuff_reg[15][12]  ( .D(n638), .CK(clk), .RN(n21), .Q(
        \gbuff[15][12] ) );
  DFFRX1 \gbuff_reg[15][11]  ( .D(n637), .CK(clk), .RN(n17), .Q(
        \gbuff[15][11] ) );
  DFFRX1 \gbuff_reg[15][10]  ( .D(n636), .CK(clk), .RN(n17), .Q(
        \gbuff[15][10] ) );
  DFFRX1 \gbuff_reg[15][9]  ( .D(n635), .CK(clk), .RN(n21), .Q(\gbuff[15][9] )
         );
  DFFRX1 \gbuff_reg[15][8]  ( .D(n634), .CK(clk), .RN(n17), .Q(\gbuff[15][8] )
         );
  DFFRX1 \gbuff_reg[15][7]  ( .D(n633), .CK(clk), .RN(n23), .Q(\gbuff[15][7] )
         );
  DFFRX1 \gbuff_reg[15][6]  ( .D(n632), .CK(clk), .RN(n24), .Q(\gbuff[15][6] )
         );
  DFFRX1 \gbuff_reg[15][5]  ( .D(n631), .CK(clk), .RN(n24), .Q(\gbuff[15][5] )
         );
  DFFRX1 \gbuff_reg[15][4]  ( .D(n630), .CK(clk), .RN(n21), .Q(\gbuff[15][4] )
         );
  DFFRX1 \gbuff_reg[15][3]  ( .D(n629), .CK(clk), .RN(n17), .Q(\gbuff[15][3] )
         );
  DFFRX1 \gbuff_reg[15][2]  ( .D(n628), .CK(clk), .RN(n24), .Q(\gbuff[15][2] )
         );
  DFFRX1 \gbuff_reg[15][1]  ( .D(n627), .CK(clk), .RN(n19), .Q(\gbuff[15][1] )
         );
  DFFRX1 \gbuff_reg[15][0]  ( .D(n626), .CK(clk), .RN(n17), .Q(\gbuff[15][0] )
         );
  DFFRX1 \gbuff_reg[11][31]  ( .D(n529), .CK(clk), .RN(n24), .Q(
        \gbuff[11][31] ) );
  DFFRX1 \gbuff_reg[11][30]  ( .D(n528), .CK(clk), .RN(n25), .Q(
        \gbuff[11][30] ) );
  DFFRX1 \gbuff_reg[11][29]  ( .D(n527), .CK(clk), .RN(n24), .Q(
        \gbuff[11][29] ) );
  DFFRX1 \gbuff_reg[11][28]  ( .D(n526), .CK(clk), .RN(n25), .Q(
        \gbuff[11][28] ) );
  DFFRX1 \gbuff_reg[11][27]  ( .D(n525), .CK(clk), .RN(n19), .Q(
        \gbuff[11][27] ) );
  DFFRX1 \gbuff_reg[11][26]  ( .D(n524), .CK(clk), .RN(n25), .Q(
        \gbuff[11][26] ) );
  DFFRX1 \gbuff_reg[11][25]  ( .D(n523), .CK(clk), .RN(n19), .Q(
        \gbuff[11][25] ) );
  DFFRX1 \gbuff_reg[11][24]  ( .D(n522), .CK(clk), .RN(n19), .Q(
        \gbuff[11][24] ) );
  DFFRX1 \gbuff_reg[11][23]  ( .D(n521), .CK(clk), .RN(n24), .Q(
        \gbuff[11][23] ) );
  DFFRX1 \gbuff_reg[11][22]  ( .D(n520), .CK(clk), .RN(n25), .Q(
        \gbuff[11][22] ) );
  DFFRX1 \gbuff_reg[11][21]  ( .D(n519), .CK(clk), .RN(n20), .Q(
        \gbuff[11][21] ) );
  DFFRX1 \gbuff_reg[11][20]  ( .D(n518), .CK(clk), .RN(n20), .Q(
        \gbuff[11][20] ) );
  DFFRX1 \gbuff_reg[11][19]  ( .D(n517), .CK(clk), .RN(n26), .Q(
        \gbuff[11][19] ) );
  DFFRX1 \gbuff_reg[11][18]  ( .D(n516), .CK(clk), .RN(n26), .Q(
        \gbuff[11][18] ) );
  DFFRX1 \gbuff_reg[11][17]  ( .D(n515), .CK(clk), .RN(n17), .Q(
        \gbuff[11][17] ) );
  DFFRX1 \gbuff_reg[11][16]  ( .D(n514), .CK(clk), .RN(n18), .Q(
        \gbuff[11][16] ) );
  DFFRX1 \gbuff_reg[11][15]  ( .D(n513), .CK(clk), .RN(n21), .Q(
        \gbuff[11][15] ) );
  DFFRX1 \gbuff_reg[11][14]  ( .D(n512), .CK(clk), .RN(n17), .Q(
        \gbuff[11][14] ) );
  DFFRX1 \gbuff_reg[11][13]  ( .D(n511), .CK(clk), .RN(n17), .Q(
        \gbuff[11][13] ) );
  DFFRX1 \gbuff_reg[11][12]  ( .D(n510), .CK(clk), .RN(n20), .Q(
        \gbuff[11][12] ) );
  DFFRX1 \gbuff_reg[11][11]  ( .D(n509), .CK(clk), .RN(n26), .Q(
        \gbuff[11][11] ) );
  DFFRX1 \gbuff_reg[11][10]  ( .D(n508), .CK(clk), .RN(n26), .Q(
        \gbuff[11][10] ) );
  DFFRX1 \gbuff_reg[11][9]  ( .D(n507), .CK(clk), .RN(n21), .Q(\gbuff[11][9] )
         );
  DFFRX1 \gbuff_reg[11][8]  ( .D(n506), .CK(clk), .RN(n18), .Q(\gbuff[11][8] )
         );
  DFFRX1 \gbuff_reg[11][7]  ( .D(n505), .CK(clk), .RN(n25), .Q(\gbuff[11][7] )
         );
  DFFRX1 \gbuff_reg[11][6]  ( .D(n504), .CK(clk), .RN(n26), .Q(\gbuff[11][6] )
         );
  DFFRX1 \gbuff_reg[11][5]  ( .D(n503), .CK(clk), .RN(n17), .Q(\gbuff[11][5] )
         );
  DFFRX1 \gbuff_reg[11][4]  ( .D(n502), .CK(clk), .RN(n23), .Q(\gbuff[11][4] )
         );
  DFFRX1 \gbuff_reg[11][3]  ( .D(n501), .CK(clk), .RN(n20), .Q(\gbuff[11][3] )
         );
  DFFRX1 \gbuff_reg[11][2]  ( .D(n500), .CK(clk), .RN(n17), .Q(\gbuff[11][2] )
         );
  DFFRX1 \gbuff_reg[11][1]  ( .D(n499), .CK(clk), .RN(n25), .Q(\gbuff[11][1] )
         );
  DFFRX1 \gbuff_reg[11][0]  ( .D(n498), .CK(clk), .RN(n23), .Q(\gbuff[11][0] )
         );
  DFFRX1 \gbuff_reg[7][31]  ( .D(n401), .CK(clk), .RN(n25), .Q(\gbuff[7][31] )
         );
  DFFRX1 \gbuff_reg[7][30]  ( .D(n400), .CK(clk), .RN(n26), .Q(\gbuff[7][30] )
         );
  DFFRX1 \gbuff_reg[7][29]  ( .D(n399), .CK(clk), .RN(n21), .Q(\gbuff[7][29] )
         );
  DFFRX1 \gbuff_reg[7][28]  ( .D(n398), .CK(clk), .RN(n19), .Q(\gbuff[7][28] )
         );
  DFFRX1 \gbuff_reg[7][27]  ( .D(n397), .CK(clk), .RN(n23), .Q(\gbuff[7][27] )
         );
  DFFRX1 \gbuff_reg[7][26]  ( .D(n396), .CK(clk), .RN(n18), .Q(\gbuff[7][26] )
         );
  DFFRX1 \gbuff_reg[7][25]  ( .D(n395), .CK(clk), .RN(n19), .Q(\gbuff[7][25] )
         );
  DFFRX1 \gbuff_reg[7][24]  ( .D(n394), .CK(clk), .RN(n20), .Q(\gbuff[7][24] )
         );
  DFFRX1 \gbuff_reg[7][23]  ( .D(n393), .CK(clk), .RN(n18), .Q(\gbuff[7][23] )
         );
  DFFRX1 \gbuff_reg[7][22]  ( .D(n392), .CK(clk), .RN(n18), .Q(\gbuff[7][22] )
         );
  DFFRX1 \gbuff_reg[7][21]  ( .D(n391), .CK(clk), .RN(n18), .Q(\gbuff[7][21] )
         );
  DFFRX1 \gbuff_reg[7][20]  ( .D(n390), .CK(clk), .RN(n18), .Q(\gbuff[7][20] )
         );
  DFFRX1 \gbuff_reg[7][19]  ( .D(n389), .CK(clk), .RN(n23), .Q(\gbuff[7][19] )
         );
  DFFRX1 \gbuff_reg[7][18]  ( .D(n388), .CK(clk), .RN(n25), .Q(\gbuff[7][18] )
         );
  DFFRX1 \gbuff_reg[7][17]  ( .D(n387), .CK(clk), .RN(n20), .Q(\gbuff[7][17] )
         );
  DFFRX1 \gbuff_reg[7][16]  ( .D(n386), .CK(clk), .RN(n20), .Q(\gbuff[7][16] )
         );
  DFFRX1 \gbuff_reg[7][15]  ( .D(n385), .CK(clk), .RN(n19), .Q(\gbuff[7][15] )
         );
  DFFRX1 \gbuff_reg[7][14]  ( .D(n384), .CK(clk), .RN(n24), .Q(\gbuff[7][14] )
         );
  DFFRX1 \gbuff_reg[7][13]  ( .D(n383), .CK(clk), .RN(n18), .Q(\gbuff[7][13] )
         );
  DFFRX1 \gbuff_reg[7][12]  ( .D(n382), .CK(clk), .RN(n26), .Q(\gbuff[7][12] )
         );
  DFFRX1 \gbuff_reg[7][11]  ( .D(n381), .CK(clk), .RN(n17), .Q(\gbuff[7][11] )
         );
  DFFRX1 \gbuff_reg[7][10]  ( .D(n380), .CK(clk), .RN(n26), .Q(\gbuff[7][10] )
         );
  DFFRX1 \gbuff_reg[7][9]  ( .D(n379), .CK(clk), .RN(n23), .Q(\gbuff[7][9] )
         );
  DFFRX1 \gbuff_reg[7][8]  ( .D(n378), .CK(clk), .RN(n25), .Q(\gbuff[7][8] )
         );
  DFFRX1 \gbuff_reg[7][7]  ( .D(n377), .CK(clk), .RN(n19), .Q(\gbuff[7][7] )
         );
  DFFRX1 \gbuff_reg[7][6]  ( .D(n376), .CK(clk), .RN(n24), .Q(\gbuff[7][6] )
         );
  DFFRX1 \gbuff_reg[7][5]  ( .D(n375), .CK(clk), .RN(n19), .Q(\gbuff[7][5] )
         );
  DFFRX1 \gbuff_reg[7][4]  ( .D(n374), .CK(clk), .RN(n21), .Q(\gbuff[7][4] )
         );
  DFFRX1 \gbuff_reg[7][3]  ( .D(n373), .CK(clk), .RN(n21), .Q(\gbuff[7][3] )
         );
  DFFRX1 \gbuff_reg[7][2]  ( .D(n372), .CK(clk), .RN(n24), .Q(\gbuff[7][2] )
         );
  DFFRX1 \gbuff_reg[7][1]  ( .D(n371), .CK(clk), .RN(n18), .Q(\gbuff[7][1] )
         );
  DFFRX1 \gbuff_reg[7][0]  ( .D(n370), .CK(clk), .RN(n21), .Q(\gbuff[7][0] )
         );
  DFFRX1 \gbuff_reg[3][31]  ( .D(n273), .CK(clk), .RN(n24), .Q(\gbuff[3][31] )
         );
  DFFRX1 \gbuff_reg[3][30]  ( .D(n272), .CK(clk), .RN(n20), .Q(\gbuff[3][30] )
         );
  DFFRX1 \gbuff_reg[3][29]  ( .D(n271), .CK(clk), .RN(n20), .Q(\gbuff[3][29] )
         );
  DFFRX1 \gbuff_reg[3][28]  ( .D(n270), .CK(clk), .RN(n17), .Q(\gbuff[3][28] )
         );
  DFFRX1 \gbuff_reg[3][27]  ( .D(n269), .CK(clk), .RN(n21), .Q(\gbuff[3][27] )
         );
  DFFRX1 \gbuff_reg[3][26]  ( .D(n268), .CK(clk), .RN(n23), .Q(\gbuff[3][26] )
         );
  DFFRX1 \gbuff_reg[3][25]  ( .D(n267), .CK(clk), .RN(n18), .Q(\gbuff[3][25] )
         );
  DFFRX1 \gbuff_reg[3][24]  ( .D(n266), .CK(clk), .RN(n21), .Q(\gbuff[3][24] )
         );
  DFFRX1 \gbuff_reg[3][23]  ( .D(n265), .CK(clk), .RN(n20), .Q(\gbuff[3][23] )
         );
  DFFRX1 \gbuff_reg[3][22]  ( .D(n264), .CK(clk), .RN(n17), .Q(\gbuff[3][22] )
         );
  DFFRX1 \gbuff_reg[3][21]  ( .D(n263), .CK(clk), .RN(n20), .Q(\gbuff[3][21] )
         );
  DFFRX1 \gbuff_reg[3][20]  ( .D(n262), .CK(clk), .RN(n25), .Q(\gbuff[3][20] )
         );
  DFFRX1 \gbuff_reg[3][19]  ( .D(n261), .CK(clk), .RN(n26), .Q(\gbuff[3][19] )
         );
  DFFRX1 \gbuff_reg[3][18]  ( .D(n260), .CK(clk), .RN(n18), .Q(\gbuff[3][18] )
         );
  DFFRX1 \gbuff_reg[3][17]  ( .D(n259), .CK(clk), .RN(n26), .Q(\gbuff[3][17] )
         );
  DFFRX1 \gbuff_reg[3][16]  ( .D(n258), .CK(clk), .RN(n26), .Q(\gbuff[3][16] )
         );
  DFFRX1 \gbuff_reg[3][15]  ( .D(n257), .CK(clk), .RN(n20), .Q(\gbuff[3][15] )
         );
  DFFRX1 \gbuff_reg[3][14]  ( .D(n256), .CK(clk), .RN(n17), .Q(\gbuff[3][14] )
         );
  DFFRX1 \gbuff_reg[3][13]  ( .D(n255), .CK(clk), .RN(n23), .Q(\gbuff[3][13] )
         );
  DFFRX1 \gbuff_reg[3][12]  ( .D(n254), .CK(clk), .RN(n23), .Q(\gbuff[3][12] )
         );
  DFFRX1 \gbuff_reg[3][11]  ( .D(n253), .CK(clk), .RN(n18), .Q(\gbuff[3][11] )
         );
  DFFRX1 \gbuff_reg[3][10]  ( .D(n252), .CK(clk), .RN(n20), .Q(\gbuff[3][10] )
         );
  DFFRX1 \gbuff_reg[3][9]  ( .D(n251), .CK(clk), .RN(n23), .Q(\gbuff[3][9] )
         );
  DFFRX1 \gbuff_reg[3][8]  ( .D(n250), .CK(clk), .RN(n19), .Q(\gbuff[3][8] )
         );
  DFFRX1 \gbuff_reg[3][7]  ( .D(n249), .CK(clk), .RN(n25), .Q(\gbuff[3][7] )
         );
  DFFRX1 \gbuff_reg[3][6]  ( .D(n248), .CK(clk), .RN(n21), .Q(\gbuff[3][6] )
         );
  DFFRX1 \gbuff_reg[3][5]  ( .D(n247), .CK(clk), .RN(n21), .Q(\gbuff[3][5] )
         );
  DFFRX1 \gbuff_reg[3][4]  ( .D(n246), .CK(clk), .RN(n24), .Q(\gbuff[3][4] )
         );
  DFFRX1 \gbuff_reg[3][3]  ( .D(n245), .CK(clk), .RN(n18), .Q(\gbuff[3][3] )
         );
  DFFRX1 \gbuff_reg[3][2]  ( .D(n244), .CK(clk), .RN(n19), .Q(\gbuff[3][2] )
         );
  DFFRX1 \gbuff_reg[3][1]  ( .D(n243), .CK(clk), .RN(n17), .Q(\gbuff[3][1] )
         );
  DFFRX1 \gbuff_reg[3][0]  ( .D(n242), .CK(clk), .RN(n19), .Q(\gbuff[3][0] )
         );
  EDFFX2 \data_out_reg[31]  ( .D(N16), .E(N81), .CK(clk), .Q(data_out[31]) );
  EDFFX2 \data_out_reg[30]  ( .D(N17), .E(N81), .CK(clk), .Q(data_out[30]) );
  EDFFX2 \data_out_reg[29]  ( .D(N18), .E(N81), .CK(clk), .Q(data_out[29]) );
  EDFFX2 \data_out_reg[28]  ( .D(N19), .E(N81), .CK(clk), .Q(data_out[28]) );
  EDFFX2 \data_out_reg[27]  ( .D(N20), .E(N81), .CK(clk), .Q(data_out[27]) );
  EDFFX2 \data_out_reg[26]  ( .D(N21), .E(N81), .CK(clk), .Q(data_out[26]) );
  EDFFX2 \data_out_reg[25]  ( .D(N22), .E(N81), .CK(clk), .Q(data_out[25]) );
  EDFFX2 \data_out_reg[24]  ( .D(N23), .E(N81), .CK(clk), .Q(data_out[24]) );
  EDFFX2 \data_out_reg[7]  ( .D(N40), .E(N81), .CK(clk), .Q(data_out[7]) );
  EDFFX2 \data_out_reg[6]  ( .D(N41), .E(N81), .CK(clk), .Q(data_out[6]) );
  EDFFX2 \data_out_reg[5]  ( .D(N42), .E(N81), .CK(clk), .Q(data_out[5]) );
  EDFFX2 \data_out_reg[4]  ( .D(N43), .E(N81), .CK(clk), .Q(data_out[4]) );
  EDFFX2 \data_out_reg[3]  ( .D(N44), .E(N81), .CK(clk), .Q(data_out[3]) );
  EDFFX2 \data_out_reg[2]  ( .D(N45), .E(N81), .CK(clk), .Q(data_out[2]) );
  EDFFX2 \data_out_reg[1]  ( .D(N46), .E(N81), .CK(clk), .Q(data_out[1]) );
  EDFFX2 \data_out_reg[0]  ( .D(N47), .E(N81), .CK(clk), .Q(data_out[0]) );
  EDFFX1 \data_out_reg[23]  ( .D(N24), .E(N81), .CK(clk), .Q(data_out[23]) );
  EDFFX1 \data_out_reg[22]  ( .D(N25), .E(N81), .CK(clk), .Q(data_out[22]) );
  EDFFX1 \data_out_reg[21]  ( .D(N26), .E(N81), .CK(clk), .Q(data_out[21]) );
  EDFFX1 \data_out_reg[20]  ( .D(N27), .E(N81), .CK(clk), .Q(data_out[20]) );
  EDFFX1 \data_out_reg[19]  ( .D(N28), .E(N81), .CK(clk), .Q(data_out[19]) );
  EDFFX1 \data_out_reg[18]  ( .D(N29), .E(N81), .CK(clk), .Q(data_out[18]) );
  EDFFX1 \data_out_reg[17]  ( .D(N30), .E(N81), .CK(clk), .Q(data_out[17]) );
  EDFFX1 \data_out_reg[16]  ( .D(N31), .E(N81), .CK(clk), .Q(data_out[16]) );
  EDFFX1 \data_out_reg[15]  ( .D(N32), .E(N81), .CK(clk), .Q(data_out[15]) );
  EDFFX1 \data_out_reg[14]  ( .D(N33), .E(N81), .CK(clk), .Q(data_out[14]) );
  EDFFX1 \data_out_reg[13]  ( .D(N34), .E(N81), .CK(clk), .Q(data_out[13]) );
  EDFFX1 \data_out_reg[12]  ( .D(N35), .E(N81), .CK(clk), .Q(data_out[12]) );
  EDFFX1 \data_out_reg[11]  ( .D(N36), .E(N81), .CK(clk), .Q(data_out[11]) );
  EDFFX1 \data_out_reg[10]  ( .D(N37), .E(N81), .CK(clk), .Q(data_out[10]) );
  EDFFX1 \data_out_reg[9]  ( .D(N38), .E(N81), .CK(clk), .Q(data_out[9]) );
  EDFFX1 \data_out_reg[8]  ( .D(N39), .E(N81), .CK(clk), .Q(data_out[8]) );
  NOR4BX1 U2 ( .AN(wr_en), .B(index[5]), .C(index[7]), .D(index[6]), .Y(n118)
         );
  NOR3BX2 U3 ( .AN(n118), .B(N13), .C(N14), .Y(n103) );
  NOR3BX2 U4 ( .AN(n118), .B(N14), .C(n1614), .Y(n120) );
  NAND2X1 U5 ( .A(n102), .B(n103), .Y(n1) );
  NAND2X1 U6 ( .A(n105), .B(n103), .Y(n2) );
  NAND2X1 U7 ( .A(n107), .B(n103), .Y(n3) );
  NAND2X1 U8 ( .A(n109), .B(n103), .Y(n4) );
  NAND2X1 U9 ( .A(n111), .B(n103), .Y(n5) );
  NAND2X1 U10 ( .A(n113), .B(n103), .Y(n6) );
  NAND2X1 U11 ( .A(n115), .B(n103), .Y(n7) );
  NAND2X1 U12 ( .A(n117), .B(n103), .Y(n8) );
  NAND2X1 U13 ( .A(n120), .B(n102), .Y(n9) );
  NAND2X1 U14 ( .A(n120), .B(n105), .Y(n10) );
  NAND2X1 U15 ( .A(n120), .B(n107), .Y(n11) );
  NAND2X1 U16 ( .A(n120), .B(n109), .Y(n12) );
  NAND2X1 U17 ( .A(n120), .B(n111), .Y(n13) );
  NAND2X1 U18 ( .A(n120), .B(n113), .Y(n14) );
  NAND2X1 U19 ( .A(n120), .B(n115), .Y(n15) );
  NAND2X1 U20 ( .A(n120), .B(n117), .Y(n16) );
  NOR2X6 U21 ( .A(wr_en), .B(rst), .Y(N81) );
  INVX20 U22 ( .A(n22), .Y(n19) );
  INVX20 U23 ( .A(n22), .Y(n21) );
  INVX20 U24 ( .A(n22), .Y(n20) );
  INVX20 U25 ( .A(n22), .Y(n17) );
  INVX20 U26 ( .A(n22), .Y(n18) );
  INVX20 U27 ( .A(n22), .Y(n25) );
  INVX20 U28 ( .A(n22), .Y(n26) );
  INVX20 U29 ( .A(n22), .Y(n24) );
  INVX20 U30 ( .A(n22), .Y(n23) );
  INVX6 U31 ( .A(n27), .Y(n22) );
  INVXL U32 ( .A(rst), .Y(n27) );
  CLKINVX1 U33 ( .A(n1610), .Y(n1609) );
  CLKINVX1 U34 ( .A(n1612), .Y(n1611) );
  CLKINVX1 U35 ( .A(N11), .Y(n1612) );
  CLKINVX1 U36 ( .A(N10), .Y(n1610) );
  CLKINVX1 U37 ( .A(N13), .Y(n1614) );
  CLKINVX1 U38 ( .A(data_in[0]), .Y(n1646) );
  CLKINVX1 U39 ( .A(data_in[1]), .Y(n1645) );
  CLKINVX1 U40 ( .A(data_in[2]), .Y(n1644) );
  CLKINVX1 U41 ( .A(data_in[3]), .Y(n1643) );
  CLKINVX1 U42 ( .A(data_in[4]), .Y(n1642) );
  CLKINVX1 U43 ( .A(data_in[5]), .Y(n1641) );
  CLKINVX1 U44 ( .A(data_in[6]), .Y(n1640) );
  CLKINVX1 U45 ( .A(data_in[7]), .Y(n1639) );
  CLKINVX1 U46 ( .A(data_in[8]), .Y(n1638) );
  CLKINVX1 U47 ( .A(data_in[9]), .Y(n1637) );
  CLKINVX1 U48 ( .A(data_in[10]), .Y(n1636) );
  CLKINVX1 U49 ( .A(data_in[11]), .Y(n1635) );
  CLKINVX1 U50 ( .A(data_in[12]), .Y(n1634) );
  CLKINVX1 U51 ( .A(data_in[13]), .Y(n1633) );
  CLKINVX1 U52 ( .A(data_in[14]), .Y(n1632) );
  CLKINVX1 U53 ( .A(data_in[15]), .Y(n1631) );
  CLKINVX1 U54 ( .A(data_in[16]), .Y(n1630) );
  CLKINVX1 U55 ( .A(data_in[17]), .Y(n1629) );
  CLKINVX1 U56 ( .A(data_in[18]), .Y(n1628) );
  CLKINVX1 U57 ( .A(data_in[19]), .Y(n1627) );
  CLKINVX1 U58 ( .A(data_in[20]), .Y(n1626) );
  CLKINVX1 U59 ( .A(data_in[21]), .Y(n1625) );
  CLKINVX1 U60 ( .A(data_in[22]), .Y(n1624) );
  CLKINVX1 U61 ( .A(data_in[23]), .Y(n1623) );
  CLKINVX1 U62 ( .A(data_in[24]), .Y(n1622) );
  CLKINVX1 U63 ( .A(data_in[25]), .Y(n1621) );
  CLKINVX1 U64 ( .A(data_in[26]), .Y(n1620) );
  CLKINVX1 U65 ( .A(data_in[27]), .Y(n1619) );
  CLKINVX1 U66 ( .A(data_in[28]), .Y(n1618) );
  CLKINVX1 U67 ( .A(data_in[29]), .Y(n1617) );
  CLKINVX1 U68 ( .A(data_in[30]), .Y(n1616) );
  CLKINVX1 U69 ( .A(data_in[31]), .Y(n1615) );
  CLKBUFX3 U70 ( .A(n1430), .Y(n1433) );
  CLKBUFX3 U71 ( .A(n1430), .Y(n1434) );
  CLKBUFX3 U72 ( .A(n1429), .Y(n1435) );
  CLKBUFX3 U73 ( .A(n1429), .Y(n1436) );
  CLKBUFX3 U74 ( .A(n1429), .Y(n1437) );
  CLKBUFX3 U75 ( .A(n1429), .Y(n1438) );
  CLKBUFX3 U76 ( .A(n1429), .Y(n1439) );
  CLKBUFX3 U77 ( .A(n1429), .Y(n1440) );
  CLKBUFX3 U78 ( .A(n1429), .Y(n1441) );
  CLKBUFX3 U79 ( .A(n1430), .Y(n1442) );
  CLKBUFX3 U80 ( .A(n1429), .Y(n1443) );
  CLKBUFX3 U81 ( .A(n1429), .Y(n1444) );
  CLKBUFX3 U82 ( .A(n1430), .Y(n1445) );
  CLKBUFX3 U83 ( .A(n1430), .Y(n1446) );
  CLKBUFX3 U84 ( .A(n1429), .Y(n1447) );
  CLKBUFX3 U85 ( .A(N11), .Y(n1412) );
  CLKBUFX3 U86 ( .A(n1410), .Y(n1413) );
  CLKBUFX3 U87 ( .A(n1410), .Y(n1414) );
  CLKBUFX3 U88 ( .A(n1410), .Y(n1415) );
  CLKBUFX3 U89 ( .A(n1410), .Y(n1416) );
  CLKBUFX3 U90 ( .A(n1410), .Y(n1417) );
  CLKBUFX3 U91 ( .A(n1410), .Y(n1418) );
  CLKBUFX3 U92 ( .A(n1410), .Y(n1419) );
  CLKBUFX3 U93 ( .A(n1410), .Y(n1420) );
  CLKBUFX3 U94 ( .A(n1410), .Y(n1421) );
  CLKBUFX3 U95 ( .A(n1410), .Y(n1422) );
  CLKBUFX3 U96 ( .A(n1410), .Y(n1423) );
  CLKBUFX3 U97 ( .A(n1611), .Y(n1424) );
  CLKBUFX3 U98 ( .A(n1410), .Y(n1425) );
  CLKBUFX3 U99 ( .A(n1410), .Y(n1426) );
  CLKBUFX3 U100 ( .A(N11), .Y(n1427) );
  CLKBUFX3 U101 ( .A(N11), .Y(n1428) );
  CLKBUFX3 U102 ( .A(n1430), .Y(n1432) );
  CLKBUFX3 U103 ( .A(n1430), .Y(n1431) );
  CLKBUFX3 U104 ( .A(N11), .Y(n1411) );
  CLKBUFX3 U105 ( .A(n1448), .Y(n1429) );
  CLKBUFX3 U106 ( .A(n1611), .Y(n1410) );
  CLKBUFX3 U107 ( .A(n1448), .Y(n1430) );
  CLKBUFX3 U108 ( .A(n1403), .Y(n1404) );
  CLKBUFX3 U109 ( .A(N13), .Y(n1405) );
  CLKBUFX3 U110 ( .A(n1403), .Y(n1406) );
  CLKBUFX3 U111 ( .A(n1613), .Y(n1407) );
  CLKBUFX3 U112 ( .A(n1613), .Y(n1408) );
  CLKBUFX3 U113 ( .A(n1613), .Y(n1409) );
  CLKBUFX3 U114 ( .A(n1609), .Y(n1448) );
  CLKBUFX3 U115 ( .A(N13), .Y(n1403) );
  CLKBUFX3 U116 ( .A(n1), .Y(n1608) );
  CLKBUFX3 U117 ( .A(n1), .Y(n1607) );
  CLKBUFX3 U118 ( .A(n2), .Y(n1604) );
  CLKBUFX3 U119 ( .A(n3), .Y(n1601) );
  CLKBUFX3 U120 ( .A(n4), .Y(n1598) );
  CLKBUFX3 U121 ( .A(n5), .Y(n1595) );
  CLKBUFX3 U122 ( .A(n6), .Y(n1592) );
  CLKBUFX3 U123 ( .A(n7), .Y(n1589) );
  CLKBUFX3 U124 ( .A(n8), .Y(n1586) );
  CLKBUFX3 U125 ( .A(n9), .Y(n1583) );
  CLKBUFX3 U126 ( .A(n10), .Y(n1580) );
  CLKBUFX3 U127 ( .A(n11), .Y(n1577) );
  CLKBUFX3 U128 ( .A(n12), .Y(n1574) );
  CLKBUFX3 U129 ( .A(n13), .Y(n1571) );
  CLKBUFX3 U130 ( .A(n14), .Y(n1568) );
  CLKBUFX3 U131 ( .A(n15), .Y(n1565) );
  CLKBUFX3 U132 ( .A(n16), .Y(n1562) );
  CLKBUFX3 U133 ( .A(n128), .Y(n1559) );
  CLKBUFX3 U134 ( .A(n130), .Y(n1556) );
  CLKBUFX3 U135 ( .A(n131), .Y(n1553) );
  CLKBUFX3 U136 ( .A(n132), .Y(n1550) );
  CLKBUFX3 U137 ( .A(n134), .Y(n1544) );
  CLKBUFX3 U138 ( .A(n135), .Y(n1541) );
  CLKBUFX3 U139 ( .A(n136), .Y(n1538) );
  CLKBUFX3 U140 ( .A(n137), .Y(n1535) );
  CLKBUFX3 U141 ( .A(n139), .Y(n1532) );
  CLKBUFX3 U142 ( .A(n140), .Y(n1529) );
  CLKBUFX3 U143 ( .A(n141), .Y(n1526) );
  CLKBUFX3 U144 ( .A(n143), .Y(n1520) );
  CLKBUFX3 U145 ( .A(n144), .Y(n1517) );
  CLKBUFX3 U146 ( .A(n145), .Y(n1514) );
  CLKBUFX3 U147 ( .A(n1), .Y(n1606) );
  CLKBUFX3 U148 ( .A(n2), .Y(n1605) );
  CLKBUFX3 U149 ( .A(n3), .Y(n1602) );
  CLKBUFX3 U150 ( .A(n4), .Y(n1599) );
  CLKBUFX3 U151 ( .A(n5), .Y(n1596) );
  CLKBUFX3 U152 ( .A(n6), .Y(n1593) );
  CLKBUFX3 U153 ( .A(n7), .Y(n1590) );
  CLKBUFX3 U154 ( .A(n8), .Y(n1587) );
  CLKBUFX3 U155 ( .A(n9), .Y(n1584) );
  CLKBUFX3 U156 ( .A(n10), .Y(n1581) );
  CLKBUFX3 U157 ( .A(n11), .Y(n1578) );
  CLKBUFX3 U158 ( .A(n12), .Y(n1575) );
  CLKBUFX3 U159 ( .A(n13), .Y(n1572) );
  CLKBUFX3 U160 ( .A(n14), .Y(n1569) );
  CLKBUFX3 U161 ( .A(n15), .Y(n1566) );
  CLKBUFX3 U162 ( .A(n16), .Y(n1563) );
  CLKBUFX3 U163 ( .A(n128), .Y(n1560) );
  CLKBUFX3 U164 ( .A(n130), .Y(n1557) );
  CLKBUFX3 U165 ( .A(n131), .Y(n1554) );
  CLKBUFX3 U166 ( .A(n132), .Y(n1551) );
  CLKBUFX3 U167 ( .A(n133), .Y(n1548) );
  CLKBUFX3 U168 ( .A(n134), .Y(n1545) );
  CLKBUFX3 U169 ( .A(n135), .Y(n1542) );
  CLKBUFX3 U170 ( .A(n136), .Y(n1539) );
  CLKBUFX3 U171 ( .A(n137), .Y(n1536) );
  CLKBUFX3 U172 ( .A(n139), .Y(n1533) );
  CLKBUFX3 U173 ( .A(n140), .Y(n1530) );
  CLKBUFX3 U174 ( .A(n141), .Y(n1527) );
  CLKBUFX3 U175 ( .A(n142), .Y(n1524) );
  CLKBUFX3 U176 ( .A(n143), .Y(n1521) );
  CLKBUFX3 U177 ( .A(n144), .Y(n1518) );
  CLKBUFX3 U178 ( .A(n145), .Y(n1515) );
  CLKBUFX3 U179 ( .A(n2), .Y(n1603) );
  CLKBUFX3 U180 ( .A(n3), .Y(n1600) );
  CLKBUFX3 U181 ( .A(n4), .Y(n1597) );
  CLKBUFX3 U182 ( .A(n5), .Y(n1594) );
  CLKBUFX3 U183 ( .A(n6), .Y(n1591) );
  CLKBUFX3 U184 ( .A(n7), .Y(n1588) );
  CLKBUFX3 U185 ( .A(n8), .Y(n1585) );
  CLKBUFX3 U186 ( .A(n9), .Y(n1582) );
  CLKBUFX3 U187 ( .A(n10), .Y(n1579) );
  CLKBUFX3 U188 ( .A(n11), .Y(n1576) );
  CLKBUFX3 U189 ( .A(n12), .Y(n1573) );
  CLKBUFX3 U190 ( .A(n13), .Y(n1570) );
  CLKBUFX3 U191 ( .A(n14), .Y(n1567) );
  CLKBUFX3 U192 ( .A(n15), .Y(n1564) );
  CLKBUFX3 U193 ( .A(n16), .Y(n1561) );
  CLKBUFX3 U194 ( .A(n128), .Y(n1558) );
  CLKBUFX3 U195 ( .A(n130), .Y(n1555) );
  CLKBUFX3 U196 ( .A(n131), .Y(n1552) );
  CLKBUFX3 U197 ( .A(n132), .Y(n1549) );
  CLKBUFX3 U198 ( .A(n133), .Y(n1546) );
  CLKBUFX3 U199 ( .A(n133), .Y(n1547) );
  CLKBUFX3 U200 ( .A(n134), .Y(n1543) );
  CLKBUFX3 U201 ( .A(n135), .Y(n1540) );
  CLKBUFX3 U202 ( .A(n136), .Y(n1537) );
  CLKBUFX3 U203 ( .A(n137), .Y(n1534) );
  CLKBUFX3 U204 ( .A(n139), .Y(n1531) );
  CLKBUFX3 U205 ( .A(n140), .Y(n1528) );
  CLKBUFX3 U206 ( .A(n141), .Y(n1525) );
  CLKBUFX3 U207 ( .A(n142), .Y(n1522) );
  CLKBUFX3 U208 ( .A(n142), .Y(n1523) );
  CLKBUFX3 U209 ( .A(n143), .Y(n1519) );
  CLKBUFX3 U210 ( .A(n144), .Y(n1516) );
  CLKBUFX3 U211 ( .A(n145), .Y(n1513) );
  CLKBUFX3 U212 ( .A(N14), .Y(n1401) );
  CLKBUFX3 U213 ( .A(N14), .Y(n1402) );
  NOR3X1 U214 ( .A(n1611), .B(n1613), .C(n1609), .Y(n102) );
  NOR3X1 U215 ( .A(n1611), .B(n1613), .C(n1610), .Y(n105) );
  NOR3X1 U216 ( .A(n1609), .B(n1613), .C(n1612), .Y(n107) );
  NOR3X1 U217 ( .A(n1610), .B(n1613), .C(n1612), .Y(n109) );
  AND3X2 U218 ( .A(n1613), .B(n1610), .C(n1612), .Y(n111) );
  AND3X2 U219 ( .A(n1613), .B(n1609), .C(n1612), .Y(n113) );
  AND3X2 U220 ( .A(n1613), .B(n1611), .C(n1610), .Y(n115) );
  AND3X2 U221 ( .A(n1613), .B(n1611), .C(n1609), .Y(n117) );
  CLKBUFX3 U222 ( .A(N12), .Y(n1613) );
  NAND2X1 U223 ( .A(n129), .B(n102), .Y(n128) );
  NAND2X1 U224 ( .A(n129), .B(n105), .Y(n130) );
  NAND2X1 U225 ( .A(n129), .B(n107), .Y(n131) );
  NAND2X1 U226 ( .A(n129), .B(n109), .Y(n132) );
  NAND2X1 U227 ( .A(n138), .B(n102), .Y(n137) );
  NAND2X1 U228 ( .A(n138), .B(n105), .Y(n139) );
  NAND2X1 U229 ( .A(n138), .B(n107), .Y(n140) );
  NAND2X1 U230 ( .A(n138), .B(n109), .Y(n141) );
  NAND2X1 U231 ( .A(n129), .B(n111), .Y(n133) );
  NAND2X1 U232 ( .A(n129), .B(n113), .Y(n134) );
  NAND2X1 U233 ( .A(n129), .B(n115), .Y(n135) );
  NAND2X1 U234 ( .A(n129), .B(n117), .Y(n136) );
  NAND2X1 U235 ( .A(n138), .B(n111), .Y(n142) );
  NAND2X1 U236 ( .A(n138), .B(n113), .Y(n143) );
  NAND2X1 U237 ( .A(n138), .B(n115), .Y(n144) );
  NAND2X1 U238 ( .A(n138), .B(n117), .Y(n145) );
  AND3X2 U239 ( .A(n118), .B(n1614), .C(N14), .Y(n129) );
  AND3X2 U240 ( .A(N13), .B(n118), .C(N14), .Y(n138) );
  CLKBUFX3 U241 ( .A(n1646), .Y(n1512) );
  CLKBUFX3 U242 ( .A(n1645), .Y(n1510) );
  CLKBUFX3 U243 ( .A(n1644), .Y(n1508) );
  CLKBUFX3 U244 ( .A(n1643), .Y(n1506) );
  CLKBUFX3 U245 ( .A(n1642), .Y(n1504) );
  CLKBUFX3 U246 ( .A(n1641), .Y(n1502) );
  CLKBUFX3 U247 ( .A(n1640), .Y(n1500) );
  CLKBUFX3 U248 ( .A(n1639), .Y(n1498) );
  CLKBUFX3 U249 ( .A(n1638), .Y(n1496) );
  CLKBUFX3 U250 ( .A(n1637), .Y(n1494) );
  CLKBUFX3 U251 ( .A(n1636), .Y(n1492) );
  CLKBUFX3 U252 ( .A(n1635), .Y(n1490) );
  CLKBUFX3 U253 ( .A(n1634), .Y(n1488) );
  CLKBUFX3 U254 ( .A(n1633), .Y(n1486) );
  CLKBUFX3 U255 ( .A(n1632), .Y(n1484) );
  CLKBUFX3 U256 ( .A(n1631), .Y(n1482) );
  CLKBUFX3 U257 ( .A(n1630), .Y(n1480) );
  CLKBUFX3 U258 ( .A(n1629), .Y(n1478) );
  CLKBUFX3 U259 ( .A(n1628), .Y(n1476) );
  CLKBUFX3 U260 ( .A(n1627), .Y(n1474) );
  CLKBUFX3 U261 ( .A(n1626), .Y(n1472) );
  CLKBUFX3 U262 ( .A(n1625), .Y(n1470) );
  CLKBUFX3 U263 ( .A(n1624), .Y(n1468) );
  CLKBUFX3 U264 ( .A(n1623), .Y(n1466) );
  CLKBUFX3 U265 ( .A(n1622), .Y(n1464) );
  CLKBUFX3 U266 ( .A(n1621), .Y(n1462) );
  CLKBUFX3 U267 ( .A(n1620), .Y(n1460) );
  CLKBUFX3 U268 ( .A(n1619), .Y(n1458) );
  CLKBUFX3 U269 ( .A(n1618), .Y(n1456) );
  CLKBUFX3 U270 ( .A(n1617), .Y(n1454) );
  CLKBUFX3 U271 ( .A(n1616), .Y(n1452) );
  CLKBUFX3 U272 ( .A(n1615), .Y(n1450) );
  CLKBUFX3 U273 ( .A(n1646), .Y(n1511) );
  CLKBUFX3 U274 ( .A(n1645), .Y(n1509) );
  CLKBUFX3 U275 ( .A(n1644), .Y(n1507) );
  CLKBUFX3 U276 ( .A(n1643), .Y(n1505) );
  CLKBUFX3 U277 ( .A(n1642), .Y(n1503) );
  CLKBUFX3 U278 ( .A(n1641), .Y(n1501) );
  CLKBUFX3 U279 ( .A(n1640), .Y(n1499) );
  CLKBUFX3 U280 ( .A(n1639), .Y(n1497) );
  CLKBUFX3 U281 ( .A(n1638), .Y(n1495) );
  CLKBUFX3 U282 ( .A(n1637), .Y(n1493) );
  CLKBUFX3 U283 ( .A(n1636), .Y(n1491) );
  CLKBUFX3 U284 ( .A(n1635), .Y(n1489) );
  CLKBUFX3 U285 ( .A(n1634), .Y(n1487) );
  CLKBUFX3 U286 ( .A(n1633), .Y(n1485) );
  CLKBUFX3 U287 ( .A(n1632), .Y(n1483) );
  CLKBUFX3 U288 ( .A(n1631), .Y(n1481) );
  CLKBUFX3 U289 ( .A(n1630), .Y(n1479) );
  CLKBUFX3 U290 ( .A(n1629), .Y(n1477) );
  CLKBUFX3 U291 ( .A(n1628), .Y(n1475) );
  CLKBUFX3 U292 ( .A(n1627), .Y(n1473) );
  CLKBUFX3 U293 ( .A(n1626), .Y(n1471) );
  CLKBUFX3 U294 ( .A(n1625), .Y(n1469) );
  CLKBUFX3 U295 ( .A(n1624), .Y(n1467) );
  CLKBUFX3 U296 ( .A(n1623), .Y(n1465) );
  CLKBUFX3 U297 ( .A(n1622), .Y(n1463) );
  CLKBUFX3 U298 ( .A(n1621), .Y(n1461) );
  CLKBUFX3 U299 ( .A(n1620), .Y(n1459) );
  CLKBUFX3 U300 ( .A(n1619), .Y(n1457) );
  CLKBUFX3 U301 ( .A(n1618), .Y(n1455) );
  CLKBUFX3 U302 ( .A(n1617), .Y(n1453) );
  CLKBUFX3 U303 ( .A(n1616), .Y(n1451) );
  CLKBUFX3 U304 ( .A(n1615), .Y(n1449) );
  MX4X1 U305 ( .A(\gbuff[4][0] ), .B(\gbuff[5][0] ), .C(\gbuff[6][0] ), .D(
        \gbuff[7][0] ), .S0(n1431), .S1(n1411), .Y(n34) );
  MX4X1 U306 ( .A(\gbuff[20][0] ), .B(\gbuff[21][0] ), .C(\gbuff[22][0] ), .D(
        \gbuff[23][0] ), .S0(n1431), .S1(n1412), .Y(n30) );
  MX4X1 U307 ( .A(\gbuff[4][1] ), .B(\gbuff[5][1] ), .C(\gbuff[6][1] ), .D(
        \gbuff[7][1] ), .S0(n1432), .S1(n1411), .Y(n44) );
  MX4X1 U308 ( .A(\gbuff[20][1] ), .B(\gbuff[21][1] ), .C(\gbuff[22][1] ), .D(
        \gbuff[23][1] ), .S0(n1432), .S1(n1411), .Y(n40) );
  MX4X1 U309 ( .A(\gbuff[4][2] ), .B(\gbuff[5][2] ), .C(\gbuff[6][2] ), .D(
        \gbuff[7][2] ), .S0(n1433), .S1(n1412), .Y(n54) );
  MX4X1 U310 ( .A(\gbuff[20][2] ), .B(\gbuff[21][2] ), .C(\gbuff[22][2] ), .D(
        \gbuff[23][2] ), .S0(n1432), .S1(n1411), .Y(n50) );
  MX4X1 U311 ( .A(\gbuff[4][3] ), .B(\gbuff[5][3] ), .C(\gbuff[6][3] ), .D(
        \gbuff[7][3] ), .S0(n1433), .S1(n1412), .Y(n64) );
  MX4X1 U312 ( .A(\gbuff[20][3] ), .B(\gbuff[21][3] ), .C(\gbuff[22][3] ), .D(
        \gbuff[23][3] ), .S0(n1433), .S1(n1412), .Y(n60) );
  MX4X1 U313 ( .A(\gbuff[4][4] ), .B(\gbuff[5][4] ), .C(\gbuff[6][4] ), .D(
        \gbuff[7][4] ), .S0(n1434), .S1(n1424), .Y(n74) );
  MX4X1 U314 ( .A(\gbuff[20][4] ), .B(\gbuff[21][4] ), .C(\gbuff[22][4] ), .D(
        \gbuff[23][4] ), .S0(n1433), .S1(n1412), .Y(n70) );
  MX4X1 U315 ( .A(\gbuff[4][5] ), .B(\gbuff[5][5] ), .C(\gbuff[6][5] ), .D(
        \gbuff[7][5] ), .S0(n1434), .S1(n1425), .Y(n84) );
  MX4X1 U316 ( .A(\gbuff[20][5] ), .B(\gbuff[21][5] ), .C(\gbuff[22][5] ), .D(
        \gbuff[23][5] ), .S0(n1434), .S1(n1426), .Y(n80) );
  MX4X1 U317 ( .A(\gbuff[4][6] ), .B(\gbuff[5][6] ), .C(\gbuff[6][6] ), .D(
        \gbuff[7][6] ), .S0(n1435), .S1(n1413), .Y(n94) );
  MX4X1 U318 ( .A(\gbuff[20][6] ), .B(\gbuff[21][6] ), .C(\gbuff[22][6] ), .D(
        \gbuff[23][6] ), .S0(n1435), .S1(n1413), .Y(n90) );
  MX4X1 U319 ( .A(\gbuff[4][7] ), .B(\gbuff[5][7] ), .C(\gbuff[6][7] ), .D(
        \gbuff[7][7] ), .S0(n1436), .S1(n1414), .Y(n108) );
  MX4X1 U320 ( .A(\gbuff[20][7] ), .B(\gbuff[21][7] ), .C(\gbuff[22][7] ), .D(
        \gbuff[23][7] ), .S0(n1435), .S1(n1413), .Y(n100) );
  MX4X1 U321 ( .A(\gbuff[4][8] ), .B(\gbuff[5][8] ), .C(\gbuff[6][8] ), .D(
        \gbuff[7][8] ), .S0(n1436), .S1(n1414), .Y(n125) );
  MX4X1 U322 ( .A(\gbuff[20][8] ), .B(\gbuff[21][8] ), .C(\gbuff[22][8] ), .D(
        \gbuff[23][8] ), .S0(n1436), .S1(n1414), .Y(n121) );
  MX4X1 U323 ( .A(\gbuff[4][9] ), .B(\gbuff[5][9] ), .C(\gbuff[6][9] ), .D(
        \gbuff[7][9] ), .S0(n1437), .S1(n1415), .Y(n1177) );
  MX4X1 U324 ( .A(\gbuff[20][9] ), .B(\gbuff[21][9] ), .C(\gbuff[22][9] ), .D(
        \gbuff[23][9] ), .S0(n1437), .S1(n1415), .Y(n1173) );
  MX4X1 U325 ( .A(\gbuff[4][10] ), .B(\gbuff[5][10] ), .C(\gbuff[6][10] ), .D(
        \gbuff[7][10] ), .S0(n1437), .S1(n1415), .Y(n1187) );
  MX4X1 U326 ( .A(\gbuff[20][10] ), .B(\gbuff[21][10] ), .C(\gbuff[22][10] ), 
        .D(\gbuff[23][10] ), .S0(n1437), .S1(n1415), .Y(n1183) );
  MX4X1 U327 ( .A(\gbuff[4][11] ), .B(\gbuff[5][11] ), .C(\gbuff[6][11] ), .D(
        \gbuff[7][11] ), .S0(n1438), .S1(n1416), .Y(n1197) );
  MX4X1 U328 ( .A(\gbuff[20][11] ), .B(\gbuff[21][11] ), .C(\gbuff[22][11] ), 
        .D(\gbuff[23][11] ), .S0(n1438), .S1(n1416), .Y(n1193) );
  MX4X1 U329 ( .A(\gbuff[4][12] ), .B(\gbuff[5][12] ), .C(\gbuff[6][12] ), .D(
        \gbuff[7][12] ), .S0(n1439), .S1(n1417), .Y(n1207) );
  MX4X1 U330 ( .A(\gbuff[20][12] ), .B(\gbuff[21][12] ), .C(\gbuff[22][12] ), 
        .D(\gbuff[23][12] ), .S0(n1438), .S1(n1416), .Y(n1203) );
  MX4X1 U331 ( .A(\gbuff[4][13] ), .B(\gbuff[5][13] ), .C(\gbuff[6][13] ), .D(
        \gbuff[7][13] ), .S0(n1439), .S1(n1417), .Y(n1217) );
  MX4X1 U332 ( .A(\gbuff[20][13] ), .B(\gbuff[21][13] ), .C(\gbuff[22][13] ), 
        .D(\gbuff[23][13] ), .S0(n1439), .S1(n1417), .Y(n1213) );
  MX4X1 U333 ( .A(\gbuff[4][14] ), .B(\gbuff[5][14] ), .C(\gbuff[6][14] ), .D(
        \gbuff[7][14] ), .S0(n1440), .S1(n1418), .Y(n1227) );
  MX4X1 U334 ( .A(\gbuff[20][14] ), .B(\gbuff[21][14] ), .C(\gbuff[22][14] ), 
        .D(\gbuff[23][14] ), .S0(n1440), .S1(n1418), .Y(n1223) );
  MX4X1 U335 ( .A(\gbuff[4][15] ), .B(\gbuff[5][15] ), .C(\gbuff[6][15] ), .D(
        \gbuff[7][15] ), .S0(n1441), .S1(n1419), .Y(n1237) );
  MX4X1 U336 ( .A(\gbuff[20][15] ), .B(\gbuff[21][15] ), .C(\gbuff[22][15] ), 
        .D(\gbuff[23][15] ), .S0(n1440), .S1(n1418), .Y(n1233) );
  MX4X1 U337 ( .A(\gbuff[4][16] ), .B(\gbuff[5][16] ), .C(\gbuff[6][16] ), .D(
        \gbuff[7][16] ), .S0(n1441), .S1(n1419), .Y(n1247) );
  MX4X1 U338 ( .A(\gbuff[20][16] ), .B(\gbuff[21][16] ), .C(\gbuff[22][16] ), 
        .D(\gbuff[23][16] ), .S0(n1441), .S1(n1419), .Y(n1243) );
  MX4X1 U339 ( .A(\gbuff[4][17] ), .B(\gbuff[5][17] ), .C(\gbuff[6][17] ), .D(
        \gbuff[7][17] ), .S0(n1442), .S1(n1420), .Y(n1257) );
  MX4X1 U340 ( .A(\gbuff[20][17] ), .B(\gbuff[21][17] ), .C(\gbuff[22][17] ), 
        .D(\gbuff[23][17] ), .S0(n1441), .S1(n1419), .Y(n1253) );
  MX4X1 U341 ( .A(\gbuff[4][18] ), .B(\gbuff[5][18] ), .C(\gbuff[6][18] ), .D(
        \gbuff[7][18] ), .S0(n1442), .S1(n1420), .Y(n1267) );
  MX4X1 U342 ( .A(\gbuff[20][18] ), .B(\gbuff[21][18] ), .C(\gbuff[22][18] ), 
        .D(\gbuff[23][18] ), .S0(n1442), .S1(n1420), .Y(n1263) );
  MX4X1 U343 ( .A(\gbuff[4][19] ), .B(\gbuff[5][19] ), .C(\gbuff[6][19] ), .D(
        \gbuff[7][19] ), .S0(n1443), .S1(n1421), .Y(n1277) );
  MX4X1 U344 ( .A(\gbuff[20][19] ), .B(\gbuff[21][19] ), .C(\gbuff[22][19] ), 
        .D(\gbuff[23][19] ), .S0(n1443), .S1(n1421), .Y(n1273) );
  MX4X1 U345 ( .A(\gbuff[4][20] ), .B(\gbuff[5][20] ), .C(\gbuff[6][20] ), .D(
        \gbuff[7][20] ), .S0(n1444), .S1(n1422), .Y(n1287) );
  MX4X1 U346 ( .A(\gbuff[20][20] ), .B(\gbuff[21][20] ), .C(\gbuff[22][20] ), 
        .D(\gbuff[23][20] ), .S0(n1443), .S1(n1421), .Y(n1283) );
  MX4X1 U347 ( .A(\gbuff[4][21] ), .B(\gbuff[5][21] ), .C(\gbuff[6][21] ), .D(
        \gbuff[7][21] ), .S0(n1444), .S1(n1422), .Y(n1297) );
  MX4X1 U348 ( .A(\gbuff[20][21] ), .B(\gbuff[21][21] ), .C(\gbuff[22][21] ), 
        .D(\gbuff[23][21] ), .S0(n1444), .S1(n1422), .Y(n1293) );
  MX4X1 U349 ( .A(\gbuff[4][22] ), .B(\gbuff[5][22] ), .C(\gbuff[6][22] ), .D(
        \gbuff[7][22] ), .S0(n1445), .S1(n1423), .Y(n1307) );
  MX4X1 U350 ( .A(\gbuff[20][22] ), .B(\gbuff[21][22] ), .C(\gbuff[22][22] ), 
        .D(\gbuff[23][22] ), .S0(n1445), .S1(n1423), .Y(n1303) );
  MX4X1 U351 ( .A(\gbuff[4][23] ), .B(\gbuff[5][23] ), .C(\gbuff[6][23] ), .D(
        \gbuff[7][23] ), .S0(n1445), .S1(n1423), .Y(n1317) );
  MX4X1 U352 ( .A(\gbuff[20][23] ), .B(\gbuff[21][23] ), .C(\gbuff[22][23] ), 
        .D(\gbuff[23][23] ), .S0(n1445), .S1(n1423), .Y(n1313) );
  MX4X1 U353 ( .A(\gbuff[4][24] ), .B(\gbuff[5][24] ), .C(\gbuff[6][24] ), .D(
        \gbuff[7][24] ), .S0(n1446), .S1(n1424), .Y(n1327) );
  MX4X1 U354 ( .A(\gbuff[20][24] ), .B(\gbuff[21][24] ), .C(\gbuff[22][24] ), 
        .D(\gbuff[23][24] ), .S0(n1446), .S1(n1424), .Y(n1323) );
  MX4X1 U355 ( .A(\gbuff[4][25] ), .B(\gbuff[5][25] ), .C(\gbuff[6][25] ), .D(
        \gbuff[7][25] ), .S0(n1429), .S1(n1425), .Y(n1337) );
  MX4X1 U356 ( .A(\gbuff[20][25] ), .B(\gbuff[21][25] ), .C(\gbuff[22][25] ), 
        .D(\gbuff[23][25] ), .S0(n1446), .S1(n1424), .Y(n1333) );
  MX4X1 U357 ( .A(\gbuff[4][26] ), .B(\gbuff[5][26] ), .C(\gbuff[6][26] ), .D(
        \gbuff[7][26] ), .S0(n1430), .S1(n1425), .Y(n1347) );
  MX4X1 U358 ( .A(\gbuff[20][26] ), .B(\gbuff[21][26] ), .C(\gbuff[22][26] ), 
        .D(\gbuff[23][26] ), .S0(n1448), .S1(n1425), .Y(n1343) );
  MX4X1 U359 ( .A(\gbuff[4][27] ), .B(\gbuff[5][27] ), .C(\gbuff[6][27] ), .D(
        \gbuff[7][27] ), .S0(n1447), .S1(n1426), .Y(n1357) );
  MX4X1 U360 ( .A(\gbuff[20][27] ), .B(\gbuff[21][27] ), .C(\gbuff[22][27] ), 
        .D(\gbuff[23][27] ), .S0(n1447), .S1(n1426), .Y(n1353) );
  MX4X1 U361 ( .A(\gbuff[4][28] ), .B(\gbuff[5][28] ), .C(\gbuff[6][28] ), .D(
        \gbuff[7][28] ), .S0(n1448), .S1(n1427), .Y(n1367) );
  MX4X1 U362 ( .A(\gbuff[20][28] ), .B(\gbuff[21][28] ), .C(\gbuff[22][28] ), 
        .D(\gbuff[23][28] ), .S0(n1447), .S1(n1426), .Y(n1363) );
  MX4X1 U363 ( .A(\gbuff[4][29] ), .B(\gbuff[5][29] ), .C(\gbuff[6][29] ), .D(
        \gbuff[7][29] ), .S0(n1448), .S1(n1427), .Y(n1377) );
  MX4X1 U364 ( .A(\gbuff[20][29] ), .B(\gbuff[21][29] ), .C(\gbuff[22][29] ), 
        .D(\gbuff[23][29] ), .S0(n1448), .S1(n1427), .Y(n1373) );
  MX4X1 U365 ( .A(\gbuff[4][30] ), .B(\gbuff[5][30] ), .C(\gbuff[6][30] ), .D(
        \gbuff[7][30] ), .S0(n1429), .S1(n1428), .Y(n1387) );
  MX4X1 U366 ( .A(\gbuff[20][30] ), .B(\gbuff[21][30] ), .C(\gbuff[22][30] ), 
        .D(\gbuff[23][30] ), .S0(n1448), .S1(n1427), .Y(n1383) );
  MX4X1 U367 ( .A(\gbuff[4][31] ), .B(\gbuff[5][31] ), .C(\gbuff[6][31] ), .D(
        \gbuff[7][31] ), .S0(n1430), .S1(n1428), .Y(n1397) );
  MX4X1 U368 ( .A(\gbuff[20][31] ), .B(\gbuff[21][31] ), .C(\gbuff[22][31] ), 
        .D(\gbuff[23][31] ), .S0(n1430), .S1(n1428), .Y(n1393) );
  MX4X1 U369 ( .A(\gbuff[0][0] ), .B(\gbuff[1][0] ), .C(\gbuff[2][0] ), .D(
        \gbuff[3][0] ), .S0(n1431), .S1(n1411), .Y(n35) );
  MX4X1 U370 ( .A(\gbuff[16][0] ), .B(\gbuff[17][0] ), .C(\gbuff[18][0] ), .D(
        \gbuff[19][0] ), .S0(n1431), .S1(n1412), .Y(n31) );
  MX4X1 U371 ( .A(\gbuff[0][1] ), .B(\gbuff[1][1] ), .C(\gbuff[2][1] ), .D(
        \gbuff[3][1] ), .S0(n1432), .S1(n1411), .Y(n45) );
  MX4X1 U372 ( .A(\gbuff[16][1] ), .B(\gbuff[17][1] ), .C(\gbuff[18][1] ), .D(
        \gbuff[19][1] ), .S0(n1432), .S1(n1411), .Y(n41) );
  MX4X1 U373 ( .A(\gbuff[0][2] ), .B(\gbuff[1][2] ), .C(\gbuff[2][2] ), .D(
        \gbuff[3][2] ), .S0(n1433), .S1(n1412), .Y(n55) );
  MX4X1 U374 ( .A(\gbuff[16][2] ), .B(\gbuff[17][2] ), .C(\gbuff[18][2] ), .D(
        \gbuff[19][2] ), .S0(n1432), .S1(n1411), .Y(n51) );
  MX4X1 U375 ( .A(\gbuff[0][3] ), .B(\gbuff[1][3] ), .C(\gbuff[2][3] ), .D(
        \gbuff[3][3] ), .S0(n1433), .S1(n1412), .Y(n65) );
  MX4X1 U376 ( .A(\gbuff[16][3] ), .B(\gbuff[17][3] ), .C(\gbuff[18][3] ), .D(
        \gbuff[19][3] ), .S0(n1433), .S1(n1412), .Y(n61) );
  MX4X1 U377 ( .A(\gbuff[0][4] ), .B(\gbuff[1][4] ), .C(\gbuff[2][4] ), .D(
        \gbuff[3][4] ), .S0(n1434), .S1(n1412), .Y(n75) );
  MX4X1 U378 ( .A(\gbuff[16][4] ), .B(\gbuff[17][4] ), .C(\gbuff[18][4] ), .D(
        \gbuff[19][4] ), .S0(n1434), .S1(n1427), .Y(n71) );
  MX4X1 U379 ( .A(\gbuff[0][5] ), .B(\gbuff[1][5] ), .C(\gbuff[2][5] ), .D(
        \gbuff[3][5] ), .S0(n1434), .S1(n1428), .Y(n85) );
  MX4X1 U380 ( .A(\gbuff[16][5] ), .B(\gbuff[17][5] ), .C(\gbuff[18][5] ), .D(
        \gbuff[19][5] ), .S0(n1434), .S1(n1411), .Y(n81) );
  MX4X1 U381 ( .A(\gbuff[0][6] ), .B(\gbuff[1][6] ), .C(\gbuff[2][6] ), .D(
        \gbuff[3][6] ), .S0(n1435), .S1(n1413), .Y(n95) );
  MX4X1 U382 ( .A(\gbuff[16][6] ), .B(\gbuff[17][6] ), .C(\gbuff[18][6] ), .D(
        \gbuff[19][6] ), .S0(n1435), .S1(n1413), .Y(n91) );
  MX4X1 U383 ( .A(\gbuff[0][7] ), .B(\gbuff[1][7] ), .C(\gbuff[2][7] ), .D(
        \gbuff[3][7] ), .S0(n1436), .S1(n1414), .Y(n110) );
  MX4X1 U384 ( .A(\gbuff[16][7] ), .B(\gbuff[17][7] ), .C(\gbuff[18][7] ), .D(
        \gbuff[19][7] ), .S0(n1435), .S1(n1413), .Y(n101) );
  MX4X1 U385 ( .A(\gbuff[0][8] ), .B(\gbuff[1][8] ), .C(\gbuff[2][8] ), .D(
        \gbuff[3][8] ), .S0(n1436), .S1(n1414), .Y(n126) );
  MX4X1 U386 ( .A(\gbuff[16][8] ), .B(\gbuff[17][8] ), .C(\gbuff[18][8] ), .D(
        \gbuff[19][8] ), .S0(n1436), .S1(n1414), .Y(n122) );
  MX4X1 U387 ( .A(\gbuff[0][9] ), .B(\gbuff[1][9] ), .C(\gbuff[2][9] ), .D(
        \gbuff[3][9] ), .S0(n1437), .S1(n1415), .Y(n1178) );
  MX4X1 U388 ( .A(\gbuff[16][9] ), .B(\gbuff[17][9] ), .C(\gbuff[18][9] ), .D(
        \gbuff[19][9] ), .S0(n1437), .S1(n1415), .Y(n1174) );
  MX4X1 U389 ( .A(\gbuff[0][10] ), .B(\gbuff[1][10] ), .C(\gbuff[2][10] ), .D(
        \gbuff[3][10] ), .S0(n1438), .S1(n1416), .Y(n1188) );
  MX4X1 U390 ( .A(\gbuff[16][10] ), .B(\gbuff[17][10] ), .C(\gbuff[18][10] ), 
        .D(\gbuff[19][10] ), .S0(n1437), .S1(n1415), .Y(n1184) );
  MX4X1 U391 ( .A(\gbuff[0][11] ), .B(\gbuff[1][11] ), .C(\gbuff[2][11] ), .D(
        \gbuff[3][11] ), .S0(n1438), .S1(n1416), .Y(n1198) );
  MX4X1 U392 ( .A(\gbuff[16][11] ), .B(\gbuff[17][11] ), .C(\gbuff[18][11] ), 
        .D(\gbuff[19][11] ), .S0(n1438), .S1(n1416), .Y(n1194) );
  MX4X1 U393 ( .A(\gbuff[0][12] ), .B(\gbuff[1][12] ), .C(\gbuff[2][12] ), .D(
        \gbuff[3][12] ), .S0(n1439), .S1(n1417), .Y(n1208) );
  MX4X1 U394 ( .A(\gbuff[16][12] ), .B(\gbuff[17][12] ), .C(\gbuff[18][12] ), 
        .D(\gbuff[19][12] ), .S0(n1438), .S1(n1416), .Y(n1204) );
  MX4X1 U395 ( .A(\gbuff[0][13] ), .B(\gbuff[1][13] ), .C(\gbuff[2][13] ), .D(
        \gbuff[3][13] ), .S0(n1439), .S1(n1417), .Y(n1218) );
  MX4X1 U396 ( .A(\gbuff[16][13] ), .B(\gbuff[17][13] ), .C(\gbuff[18][13] ), 
        .D(\gbuff[19][13] ), .S0(n1439), .S1(n1417), .Y(n1214) );
  MX4X1 U397 ( .A(\gbuff[0][14] ), .B(\gbuff[1][14] ), .C(\gbuff[2][14] ), .D(
        \gbuff[3][14] ), .S0(n1440), .S1(n1418), .Y(n1228) );
  MX4X1 U398 ( .A(\gbuff[16][14] ), .B(\gbuff[17][14] ), .C(\gbuff[18][14] ), 
        .D(\gbuff[19][14] ), .S0(n1440), .S1(n1418), .Y(n1224) );
  MX4X1 U399 ( .A(\gbuff[0][15] ), .B(\gbuff[1][15] ), .C(\gbuff[2][15] ), .D(
        \gbuff[3][15] ), .S0(n1441), .S1(n1419), .Y(n1238) );
  MX4X1 U400 ( .A(\gbuff[16][15] ), .B(\gbuff[17][15] ), .C(\gbuff[18][15] ), 
        .D(\gbuff[19][15] ), .S0(n1440), .S1(n1418), .Y(n1234) );
  MX4X1 U401 ( .A(\gbuff[0][16] ), .B(\gbuff[1][16] ), .C(\gbuff[2][16] ), .D(
        \gbuff[3][16] ), .S0(n1441), .S1(n1419), .Y(n1248) );
  MX4X1 U402 ( .A(\gbuff[16][16] ), .B(\gbuff[17][16] ), .C(\gbuff[18][16] ), 
        .D(\gbuff[19][16] ), .S0(n1441), .S1(n1419), .Y(n1244) );
  MX4X1 U403 ( .A(\gbuff[0][17] ), .B(\gbuff[1][17] ), .C(\gbuff[2][17] ), .D(
        \gbuff[3][17] ), .S0(n1442), .S1(n1420), .Y(n1258) );
  MX4X1 U404 ( .A(\gbuff[16][17] ), .B(\gbuff[17][17] ), .C(\gbuff[18][17] ), 
        .D(\gbuff[19][17] ), .S0(n1442), .S1(n1420), .Y(n1254) );
  MX4X1 U405 ( .A(\gbuff[0][18] ), .B(\gbuff[1][18] ), .C(\gbuff[2][18] ), .D(
        \gbuff[3][18] ), .S0(n1442), .S1(n1420), .Y(n1268) );
  MX4X1 U406 ( .A(\gbuff[16][18] ), .B(\gbuff[17][18] ), .C(\gbuff[18][18] ), 
        .D(\gbuff[19][18] ), .S0(n1442), .S1(n1420), .Y(n1264) );
  MX4X1 U407 ( .A(\gbuff[0][19] ), .B(\gbuff[1][19] ), .C(\gbuff[2][19] ), .D(
        \gbuff[3][19] ), .S0(n1443), .S1(n1421), .Y(n1278) );
  MX4X1 U408 ( .A(\gbuff[16][19] ), .B(\gbuff[17][19] ), .C(\gbuff[18][19] ), 
        .D(\gbuff[19][19] ), .S0(n1443), .S1(n1421), .Y(n1274) );
  MX4X1 U409 ( .A(\gbuff[0][20] ), .B(\gbuff[1][20] ), .C(\gbuff[2][20] ), .D(
        \gbuff[3][20] ), .S0(n1444), .S1(n1422), .Y(n1288) );
  MX4X1 U410 ( .A(\gbuff[16][20] ), .B(\gbuff[17][20] ), .C(\gbuff[18][20] ), 
        .D(\gbuff[19][20] ), .S0(n1443), .S1(n1421), .Y(n1284) );
  MX4X1 U411 ( .A(\gbuff[0][21] ), .B(\gbuff[1][21] ), .C(\gbuff[2][21] ), .D(
        \gbuff[3][21] ), .S0(n1444), .S1(n1422), .Y(n1298) );
  MX4X1 U412 ( .A(\gbuff[16][21] ), .B(\gbuff[17][21] ), .C(\gbuff[18][21] ), 
        .D(\gbuff[19][21] ), .S0(n1444), .S1(n1422), .Y(n1294) );
  MX4X1 U413 ( .A(\gbuff[0][22] ), .B(\gbuff[1][22] ), .C(\gbuff[2][22] ), .D(
        \gbuff[3][22] ), .S0(n1445), .S1(n1423), .Y(n1308) );
  MX4X1 U414 ( .A(\gbuff[16][22] ), .B(\gbuff[17][22] ), .C(\gbuff[18][22] ), 
        .D(\gbuff[19][22] ), .S0(n1445), .S1(n1423), .Y(n1304) );
  MX4X1 U415 ( .A(\gbuff[0][23] ), .B(\gbuff[1][23] ), .C(\gbuff[2][23] ), .D(
        \gbuff[3][23] ), .S0(n1446), .S1(n1424), .Y(n1318) );
  MX4X1 U416 ( .A(\gbuff[16][23] ), .B(\gbuff[17][23] ), .C(\gbuff[18][23] ), 
        .D(\gbuff[19][23] ), .S0(n1445), .S1(n1423), .Y(n1314) );
  MX4X1 U417 ( .A(\gbuff[0][24] ), .B(\gbuff[1][24] ), .C(\gbuff[2][24] ), .D(
        \gbuff[3][24] ), .S0(n1446), .S1(n1424), .Y(n1328) );
  MX4X1 U418 ( .A(\gbuff[16][24] ), .B(\gbuff[17][24] ), .C(\gbuff[18][24] ), 
        .D(\gbuff[19][24] ), .S0(n1446), .S1(n1424), .Y(n1324) );
  MX4X1 U419 ( .A(\gbuff[0][25] ), .B(\gbuff[1][25] ), .C(\gbuff[2][25] ), .D(
        \gbuff[3][25] ), .S0(n1431), .S1(n1425), .Y(n1338) );
  MX4X1 U420 ( .A(\gbuff[16][25] ), .B(\gbuff[17][25] ), .C(\gbuff[18][25] ), 
        .D(\gbuff[19][25] ), .S0(n1446), .S1(n1424), .Y(n1334) );
  MX4X1 U421 ( .A(\gbuff[0][26] ), .B(\gbuff[1][26] ), .C(\gbuff[2][26] ), .D(
        \gbuff[3][26] ), .S0(N10), .S1(n1425), .Y(n1348) );
  MX4X1 U422 ( .A(\gbuff[16][26] ), .B(\gbuff[17][26] ), .C(\gbuff[18][26] ), 
        .D(\gbuff[19][26] ), .S0(N10), .S1(n1425), .Y(n1344) );
  MX4X1 U423 ( .A(\gbuff[0][27] ), .B(\gbuff[1][27] ), .C(\gbuff[2][27] ), .D(
        \gbuff[3][27] ), .S0(n1447), .S1(n1426), .Y(n1358) );
  MX4X1 U424 ( .A(\gbuff[16][27] ), .B(\gbuff[17][27] ), .C(\gbuff[18][27] ), 
        .D(\gbuff[19][27] ), .S0(n1447), .S1(n1426), .Y(n1354) );
  MX4X1 U425 ( .A(\gbuff[0][28] ), .B(\gbuff[1][28] ), .C(\gbuff[2][28] ), .D(
        \gbuff[3][28] ), .S0(n1448), .S1(n1427), .Y(n1368) );
  MX4X1 U426 ( .A(\gbuff[16][28] ), .B(\gbuff[17][28] ), .C(\gbuff[18][28] ), 
        .D(\gbuff[19][28] ), .S0(n1447), .S1(n1426), .Y(n1364) );
  MX4X1 U427 ( .A(\gbuff[0][29] ), .B(\gbuff[1][29] ), .C(\gbuff[2][29] ), .D(
        \gbuff[3][29] ), .S0(n1609), .S1(n1427), .Y(n1378) );
  MX4X1 U428 ( .A(\gbuff[16][29] ), .B(\gbuff[17][29] ), .C(\gbuff[18][29] ), 
        .D(\gbuff[19][29] ), .S0(n1448), .S1(n1427), .Y(n1374) );
  MX4X1 U429 ( .A(\gbuff[0][30] ), .B(\gbuff[1][30] ), .C(\gbuff[2][30] ), .D(
        \gbuff[3][30] ), .S0(n1430), .S1(n1428), .Y(n1388) );
  MX4X1 U430 ( .A(\gbuff[16][30] ), .B(\gbuff[17][30] ), .C(\gbuff[18][30] ), 
        .D(\gbuff[19][30] ), .S0(n1430), .S1(n1428), .Y(n1384) );
  MX4X1 U431 ( .A(\gbuff[0][31] ), .B(\gbuff[1][31] ), .C(\gbuff[2][31] ), .D(
        \gbuff[3][31] ), .S0(n1429), .S1(n1428), .Y(n1398) );
  MX4X1 U432 ( .A(\gbuff[16][31] ), .B(\gbuff[17][31] ), .C(\gbuff[18][31] ), 
        .D(\gbuff[19][31] ), .S0(n1429), .S1(n1428), .Y(n1394) );
  MX4X1 U433 ( .A(\gbuff[8][0] ), .B(\gbuff[9][0] ), .C(\gbuff[10][0] ), .D(
        \gbuff[11][0] ), .S0(n1431), .S1(n1427), .Y(n33) );
  MX4X1 U434 ( .A(\gbuff[24][0] ), .B(\gbuff[25][0] ), .C(\gbuff[26][0] ), .D(
        \gbuff[27][0] ), .S0(n1431), .S1(n1428), .Y(n29) );
  MX4X1 U435 ( .A(\gbuff[8][1] ), .B(\gbuff[9][1] ), .C(\gbuff[10][1] ), .D(
        \gbuff[11][1] ), .S0(n1432), .S1(n1411), .Y(n43) );
  MX4X1 U436 ( .A(\gbuff[24][1] ), .B(\gbuff[25][1] ), .C(\gbuff[26][1] ), .D(
        \gbuff[27][1] ), .S0(n1432), .S1(n1411), .Y(n39) );
  MX4X1 U437 ( .A(\gbuff[8][2] ), .B(\gbuff[9][2] ), .C(\gbuff[10][2] ), .D(
        \gbuff[11][2] ), .S0(n1432), .S1(n1411), .Y(n53) );
  MX4X1 U438 ( .A(\gbuff[24][2] ), .B(\gbuff[25][2] ), .C(\gbuff[26][2] ), .D(
        \gbuff[27][2] ), .S0(n1432), .S1(n1411), .Y(n49) );
  MX4X1 U439 ( .A(\gbuff[8][3] ), .B(\gbuff[9][3] ), .C(\gbuff[10][3] ), .D(
        \gbuff[11][3] ), .S0(n1433), .S1(n1412), .Y(n63) );
  MX4X1 U440 ( .A(\gbuff[24][3] ), .B(\gbuff[25][3] ), .C(\gbuff[26][3] ), .D(
        \gbuff[27][3] ), .S0(n1433), .S1(n1412), .Y(n59) );
  MX4X1 U441 ( .A(\gbuff[8][4] ), .B(\gbuff[9][4] ), .C(\gbuff[10][4] ), .D(
        \gbuff[11][4] ), .S0(n1434), .S1(n1428), .Y(n73) );
  MX4X1 U442 ( .A(\gbuff[24][4] ), .B(\gbuff[25][4] ), .C(\gbuff[26][4] ), .D(
        \gbuff[27][4] ), .S0(n1433), .S1(n1412), .Y(n69) );
  MX4X1 U443 ( .A(\gbuff[8][5] ), .B(\gbuff[9][5] ), .C(\gbuff[10][5] ), .D(
        \gbuff[11][5] ), .S0(n1434), .S1(n1427), .Y(n83) );
  MX4X1 U444 ( .A(\gbuff[24][5] ), .B(\gbuff[25][5] ), .C(\gbuff[26][5] ), .D(
        \gbuff[27][5] ), .S0(n1434), .S1(n1411), .Y(n79) );
  MX4X1 U445 ( .A(\gbuff[8][6] ), .B(\gbuff[9][6] ), .C(\gbuff[10][6] ), .D(
        \gbuff[11][6] ), .S0(n1435), .S1(n1413), .Y(n93) );
  MX4X1 U446 ( .A(\gbuff[24][6] ), .B(\gbuff[25][6] ), .C(\gbuff[26][6] ), .D(
        \gbuff[27][6] ), .S0(n1435), .S1(n1413), .Y(n89) );
  MX4X1 U447 ( .A(\gbuff[8][7] ), .B(\gbuff[9][7] ), .C(\gbuff[10][7] ), .D(
        \gbuff[11][7] ), .S0(n1436), .S1(n1414), .Y(n106) );
  MX4X1 U448 ( .A(\gbuff[24][7] ), .B(\gbuff[25][7] ), .C(\gbuff[26][7] ), .D(
        \gbuff[27][7] ), .S0(n1435), .S1(n1413), .Y(n99) );
  MX4X1 U449 ( .A(\gbuff[8][8] ), .B(\gbuff[9][8] ), .C(\gbuff[10][8] ), .D(
        \gbuff[11][8] ), .S0(n1436), .S1(n1414), .Y(n124) );
  MX4X1 U450 ( .A(\gbuff[24][8] ), .B(\gbuff[25][8] ), .C(\gbuff[26][8] ), .D(
        \gbuff[27][8] ), .S0(n1436), .S1(n1414), .Y(n119) );
  MX4X1 U451 ( .A(\gbuff[8][9] ), .B(\gbuff[9][9] ), .C(\gbuff[10][9] ), .D(
        \gbuff[11][9] ), .S0(n1437), .S1(n1415), .Y(n1176) );
  MX4X1 U452 ( .A(\gbuff[24][9] ), .B(\gbuff[25][9] ), .C(\gbuff[26][9] ), .D(
        \gbuff[27][9] ), .S0(n1436), .S1(n1414), .Y(n1172) );
  MX4X1 U453 ( .A(\gbuff[8][10] ), .B(\gbuff[9][10] ), .C(\gbuff[10][10] ), 
        .D(\gbuff[11][10] ), .S0(n1437), .S1(n1415), .Y(n1186) );
  MX4X1 U454 ( .A(\gbuff[24][10] ), .B(\gbuff[25][10] ), .C(\gbuff[26][10] ), 
        .D(\gbuff[27][10] ), .S0(n1437), .S1(n1415), .Y(n1182) );
  MX4X1 U455 ( .A(\gbuff[8][11] ), .B(\gbuff[9][11] ), .C(\gbuff[10][11] ), 
        .D(\gbuff[11][11] ), .S0(n1438), .S1(n1416), .Y(n1196) );
  MX4X1 U456 ( .A(\gbuff[24][11] ), .B(\gbuff[25][11] ), .C(\gbuff[26][11] ), 
        .D(\gbuff[27][11] ), .S0(n1438), .S1(n1416), .Y(n1192) );
  MX4X1 U457 ( .A(\gbuff[8][12] ), .B(\gbuff[9][12] ), .C(\gbuff[10][12] ), 
        .D(\gbuff[11][12] ), .S0(n1439), .S1(n1417), .Y(n1206) );
  MX4X1 U458 ( .A(\gbuff[24][12] ), .B(\gbuff[25][12] ), .C(\gbuff[26][12] ), 
        .D(\gbuff[27][12] ), .S0(n1438), .S1(n1416), .Y(n1202) );
  MX4X1 U459 ( .A(\gbuff[8][13] ), .B(\gbuff[9][13] ), .C(\gbuff[10][13] ), 
        .D(\gbuff[11][13] ), .S0(n1439), .S1(n1417), .Y(n1216) );
  MX4X1 U460 ( .A(\gbuff[24][13] ), .B(\gbuff[25][13] ), .C(\gbuff[26][13] ), 
        .D(\gbuff[27][13] ), .S0(n1439), .S1(n1417), .Y(n1212) );
  MX4X1 U461 ( .A(\gbuff[8][14] ), .B(\gbuff[9][14] ), .C(\gbuff[10][14] ), 
        .D(\gbuff[11][14] ), .S0(n1440), .S1(n1418), .Y(n1226) );
  MX4X1 U462 ( .A(\gbuff[24][14] ), .B(\gbuff[25][14] ), .C(\gbuff[26][14] ), 
        .D(\gbuff[27][14] ), .S0(n1440), .S1(n1418), .Y(n1222) );
  MX4X1 U463 ( .A(\gbuff[8][15] ), .B(\gbuff[9][15] ), .C(\gbuff[10][15] ), 
        .D(\gbuff[11][15] ), .S0(n1440), .S1(n1418), .Y(n1236) );
  MX4X1 U464 ( .A(\gbuff[24][15] ), .B(\gbuff[25][15] ), .C(\gbuff[26][15] ), 
        .D(\gbuff[27][15] ), .S0(n1440), .S1(n1418), .Y(n1232) );
  MX4X1 U465 ( .A(\gbuff[8][16] ), .B(\gbuff[9][16] ), .C(\gbuff[10][16] ), 
        .D(\gbuff[11][16] ), .S0(n1441), .S1(n1419), .Y(n1246) );
  MX4X1 U466 ( .A(\gbuff[24][16] ), .B(\gbuff[25][16] ), .C(\gbuff[26][16] ), 
        .D(\gbuff[27][16] ), .S0(n1441), .S1(n1419), .Y(n1242) );
  MX4X1 U467 ( .A(\gbuff[8][17] ), .B(\gbuff[9][17] ), .C(\gbuff[10][17] ), 
        .D(\gbuff[11][17] ), .S0(n1442), .S1(n1420), .Y(n1256) );
  MX4X1 U468 ( .A(\gbuff[24][17] ), .B(\gbuff[25][17] ), .C(\gbuff[26][17] ), 
        .D(\gbuff[27][17] ), .S0(n1441), .S1(n1419), .Y(n1252) );
  MX4X1 U469 ( .A(\gbuff[8][18] ), .B(\gbuff[9][18] ), .C(\gbuff[10][18] ), 
        .D(\gbuff[11][18] ), .S0(n1442), .S1(n1420), .Y(n1266) );
  MX4X1 U470 ( .A(\gbuff[24][18] ), .B(\gbuff[25][18] ), .C(\gbuff[26][18] ), 
        .D(\gbuff[27][18] ), .S0(n1442), .S1(n1420), .Y(n1262) );
  MX4X1 U471 ( .A(\gbuff[8][19] ), .B(\gbuff[9][19] ), .C(\gbuff[10][19] ), 
        .D(\gbuff[11][19] ), .S0(n1443), .S1(n1421), .Y(n1276) );
  MX4X1 U472 ( .A(\gbuff[24][19] ), .B(\gbuff[25][19] ), .C(\gbuff[26][19] ), 
        .D(\gbuff[27][19] ), .S0(n1443), .S1(n1421), .Y(n1272) );
  MX4X1 U473 ( .A(\gbuff[8][20] ), .B(\gbuff[9][20] ), .C(\gbuff[10][20] ), 
        .D(\gbuff[11][20] ), .S0(n1444), .S1(n1422), .Y(n1286) );
  MX4X1 U474 ( .A(\gbuff[24][20] ), .B(\gbuff[25][20] ), .C(\gbuff[26][20] ), 
        .D(\gbuff[27][20] ), .S0(n1443), .S1(n1421), .Y(n1282) );
  MX4X1 U475 ( .A(\gbuff[8][21] ), .B(\gbuff[9][21] ), .C(\gbuff[10][21] ), 
        .D(\gbuff[11][21] ), .S0(n1444), .S1(n1422), .Y(n1296) );
  MX4X1 U476 ( .A(\gbuff[24][21] ), .B(\gbuff[25][21] ), .C(\gbuff[26][21] ), 
        .D(\gbuff[27][21] ), .S0(n1444), .S1(n1422), .Y(n1292) );
  MX4X1 U477 ( .A(\gbuff[8][22] ), .B(\gbuff[9][22] ), .C(\gbuff[10][22] ), 
        .D(\gbuff[11][22] ), .S0(n1445), .S1(n1423), .Y(n1306) );
  MX4X1 U478 ( .A(\gbuff[24][22] ), .B(\gbuff[25][22] ), .C(\gbuff[26][22] ), 
        .D(\gbuff[27][22] ), .S0(n1444), .S1(n1422), .Y(n1302) );
  MX4X1 U479 ( .A(\gbuff[8][23] ), .B(\gbuff[9][23] ), .C(\gbuff[10][23] ), 
        .D(\gbuff[11][23] ), .S0(n1445), .S1(n1423), .Y(n1316) );
  MX4X1 U480 ( .A(\gbuff[24][23] ), .B(\gbuff[25][23] ), .C(\gbuff[26][23] ), 
        .D(\gbuff[27][23] ), .S0(n1445), .S1(n1423), .Y(n1312) );
  MX4X1 U481 ( .A(\gbuff[8][24] ), .B(\gbuff[9][24] ), .C(\gbuff[10][24] ), 
        .D(\gbuff[11][24] ), .S0(n1446), .S1(n1424), .Y(n1326) );
  MX4X1 U482 ( .A(\gbuff[24][24] ), .B(\gbuff[25][24] ), .C(\gbuff[26][24] ), 
        .D(\gbuff[27][24] ), .S0(n1446), .S1(n1424), .Y(n1322) );
  MX4X1 U483 ( .A(\gbuff[8][25] ), .B(\gbuff[9][25] ), .C(\gbuff[10][25] ), 
        .D(\gbuff[11][25] ), .S0(n1431), .S1(n1425), .Y(n1336) );
  MX4X1 U484 ( .A(\gbuff[24][25] ), .B(\gbuff[25][25] ), .C(\gbuff[26][25] ), 
        .D(\gbuff[27][25] ), .S0(n1446), .S1(n1424), .Y(n1332) );
  MX4X1 U485 ( .A(\gbuff[8][26] ), .B(\gbuff[9][26] ), .C(\gbuff[10][26] ), 
        .D(\gbuff[11][26] ), .S0(n1431), .S1(n1425), .Y(n1346) );
  MX4X1 U486 ( .A(\gbuff[24][26] ), .B(\gbuff[25][26] ), .C(\gbuff[26][26] ), 
        .D(\gbuff[27][26] ), .S0(n1431), .S1(n1425), .Y(n1342) );
  MX4X1 U487 ( .A(\gbuff[8][27] ), .B(\gbuff[9][27] ), .C(\gbuff[10][27] ), 
        .D(\gbuff[11][27] ), .S0(n1447), .S1(n1426), .Y(n1356) );
  MX4X1 U488 ( .A(\gbuff[24][27] ), .B(\gbuff[25][27] ), .C(\gbuff[26][27] ), 
        .D(\gbuff[27][27] ), .S0(n1447), .S1(n1426), .Y(n1352) );
  MX4X1 U489 ( .A(\gbuff[8][28] ), .B(\gbuff[9][28] ), .C(\gbuff[10][28] ), 
        .D(\gbuff[11][28] ), .S0(n1447), .S1(n1426), .Y(n1366) );
  MX4X1 U490 ( .A(\gbuff[24][28] ), .B(\gbuff[25][28] ), .C(\gbuff[26][28] ), 
        .D(\gbuff[27][28] ), .S0(n1447), .S1(n1426), .Y(n1362) );
  MX4X1 U491 ( .A(\gbuff[8][29] ), .B(\gbuff[9][29] ), .C(\gbuff[10][29] ), 
        .D(\gbuff[11][29] ), .S0(n1429), .S1(n1427), .Y(n1376) );
  MX4X1 U492 ( .A(\gbuff[24][29] ), .B(\gbuff[25][29] ), .C(\gbuff[26][29] ), 
        .D(\gbuff[27][29] ), .S0(n1430), .S1(n1427), .Y(n1372) );
  MX4X1 U493 ( .A(\gbuff[8][30] ), .B(\gbuff[9][30] ), .C(\gbuff[10][30] ), 
        .D(\gbuff[11][30] ), .S0(n1430), .S1(n1428), .Y(n1386) );
  MX4X1 U494 ( .A(\gbuff[24][30] ), .B(\gbuff[25][30] ), .C(\gbuff[26][30] ), 
        .D(\gbuff[27][30] ), .S0(n1448), .S1(n1427), .Y(n1382) );
  MX4X1 U495 ( .A(\gbuff[8][31] ), .B(\gbuff[9][31] ), .C(\gbuff[10][31] ), 
        .D(\gbuff[11][31] ), .S0(n1448), .S1(n1428), .Y(n1396) );
  MX4X1 U496 ( .A(\gbuff[24][31] ), .B(\gbuff[25][31] ), .C(\gbuff[26][31] ), 
        .D(\gbuff[27][31] ), .S0(n1429), .S1(n1428), .Y(n1392) );
  MX4X1 U497 ( .A(\gbuff[12][0] ), .B(\gbuff[13][0] ), .C(\gbuff[14][0] ), .D(
        \gbuff[15][0] ), .S0(n1431), .S1(n1424), .Y(n32) );
  MX4X1 U498 ( .A(\gbuff[12][1] ), .B(\gbuff[13][1] ), .C(\gbuff[14][1] ), .D(
        \gbuff[15][1] ), .S0(n1432), .S1(n1411), .Y(n42) );
  MX4X1 U499 ( .A(\gbuff[12][2] ), .B(\gbuff[13][2] ), .C(\gbuff[14][2] ), .D(
        \gbuff[15][2] ), .S0(n1432), .S1(n1411), .Y(n52) );
  MX4X1 U500 ( .A(\gbuff[12][3] ), .B(\gbuff[13][3] ), .C(\gbuff[14][3] ), .D(
        \gbuff[15][3] ), .S0(n1433), .S1(n1412), .Y(n62) );
  MX4X1 U501 ( .A(\gbuff[12][4] ), .B(\gbuff[13][4] ), .C(\gbuff[14][4] ), .D(
        \gbuff[15][4] ), .S0(n1434), .S1(n1412), .Y(n72) );
  MX4X1 U502 ( .A(\gbuff[12][5] ), .B(\gbuff[13][5] ), .C(\gbuff[14][5] ), .D(
        \gbuff[15][5] ), .S0(n1434), .S1(n1424), .Y(n82) );
  MX4X1 U503 ( .A(\gbuff[12][6] ), .B(\gbuff[13][6] ), .C(\gbuff[14][6] ), .D(
        \gbuff[15][6] ), .S0(n1435), .S1(n1413), .Y(n92) );
  MX4X1 U504 ( .A(\gbuff[12][7] ), .B(\gbuff[13][7] ), .C(\gbuff[14][7] ), .D(
        \gbuff[15][7] ), .S0(n1435), .S1(n1413), .Y(n104) );
  MX4X1 U505 ( .A(\gbuff[12][8] ), .B(\gbuff[13][8] ), .C(\gbuff[14][8] ), .D(
        \gbuff[15][8] ), .S0(n1436), .S1(n1414), .Y(n123) );
  MX4X1 U506 ( .A(\gbuff[12][9] ), .B(\gbuff[13][9] ), .C(\gbuff[14][9] ), .D(
        \gbuff[15][9] ), .S0(n1437), .S1(n1415), .Y(n1175) );
  MX4X1 U507 ( .A(\gbuff[12][10] ), .B(\gbuff[13][10] ), .C(\gbuff[14][10] ), 
        .D(\gbuff[15][10] ), .S0(n1437), .S1(n1415), .Y(n1185) );
  MX4X1 U508 ( .A(\gbuff[12][11] ), .B(\gbuff[13][11] ), .C(\gbuff[14][11] ), 
        .D(\gbuff[15][11] ), .S0(n1438), .S1(n1416), .Y(n1195) );
  MX4X1 U509 ( .A(\gbuff[12][12] ), .B(\gbuff[13][12] ), .C(\gbuff[14][12] ), 
        .D(\gbuff[15][12] ), .S0(n1439), .S1(n1417), .Y(n1205) );
  MX4X1 U510 ( .A(\gbuff[12][13] ), .B(\gbuff[13][13] ), .C(\gbuff[14][13] ), 
        .D(\gbuff[15][13] ), .S0(n1439), .S1(n1417), .Y(n1215) );
  MX4X1 U511 ( .A(\gbuff[12][14] ), .B(\gbuff[13][14] ), .C(\gbuff[14][14] ), 
        .D(\gbuff[15][14] ), .S0(n1440), .S1(n1418), .Y(n1225) );
  MX4X1 U512 ( .A(\gbuff[12][15] ), .B(\gbuff[13][15] ), .C(\gbuff[14][15] ), 
        .D(\gbuff[15][15] ), .S0(n1440), .S1(n1418), .Y(n1235) );
  MX4X1 U513 ( .A(\gbuff[12][16] ), .B(\gbuff[13][16] ), .C(\gbuff[14][16] ), 
        .D(\gbuff[15][16] ), .S0(n1441), .S1(n1419), .Y(n1245) );
  MX4X1 U514 ( .A(\gbuff[12][17] ), .B(\gbuff[13][17] ), .C(\gbuff[14][17] ), 
        .D(\gbuff[15][17] ), .S0(n1442), .S1(n1420), .Y(n1255) );
  MX4X1 U515 ( .A(\gbuff[12][18] ), .B(\gbuff[13][18] ), .C(\gbuff[14][18] ), 
        .D(\gbuff[15][18] ), .S0(n1442), .S1(n1420), .Y(n1265) );
  MX4X1 U516 ( .A(\gbuff[12][19] ), .B(\gbuff[13][19] ), .C(\gbuff[14][19] ), 
        .D(\gbuff[15][19] ), .S0(n1443), .S1(n1421), .Y(n1275) );
  MX4X1 U517 ( .A(\gbuff[12][20] ), .B(\gbuff[13][20] ), .C(\gbuff[14][20] ), 
        .D(\gbuff[15][20] ), .S0(n1443), .S1(n1421), .Y(n1285) );
  MX4X1 U518 ( .A(\gbuff[12][21] ), .B(\gbuff[13][21] ), .C(\gbuff[14][21] ), 
        .D(\gbuff[15][21] ), .S0(n1444), .S1(n1422), .Y(n1295) );
  MX4X1 U519 ( .A(\gbuff[12][22] ), .B(\gbuff[13][22] ), .C(\gbuff[14][22] ), 
        .D(\gbuff[15][22] ), .S0(n1445), .S1(n1423), .Y(n1305) );
  MX4X1 U520 ( .A(\gbuff[12][23] ), .B(\gbuff[13][23] ), .C(\gbuff[14][23] ), 
        .D(\gbuff[15][23] ), .S0(n1445), .S1(n1423), .Y(n1315) );
  MX4X1 U521 ( .A(\gbuff[12][24] ), .B(\gbuff[13][24] ), .C(\gbuff[14][24] ), 
        .D(\gbuff[15][24] ), .S0(n1446), .S1(n1424), .Y(n1325) );
  MX4X1 U522 ( .A(\gbuff[12][25] ), .B(\gbuff[13][25] ), .C(\gbuff[14][25] ), 
        .D(\gbuff[15][25] ), .S0(N10), .S1(n1425), .Y(n1335) );
  MX4X1 U523 ( .A(\gbuff[12][26] ), .B(\gbuff[13][26] ), .C(\gbuff[14][26] ), 
        .D(\gbuff[15][26] ), .S0(N10), .S1(n1425), .Y(n1345) );
  MX4X1 U524 ( .A(\gbuff[12][27] ), .B(\gbuff[13][27] ), .C(\gbuff[14][27] ), 
        .D(\gbuff[15][27] ), .S0(n1447), .S1(n1426), .Y(n1355) );
  MX4X1 U525 ( .A(\gbuff[12][28] ), .B(\gbuff[13][28] ), .C(\gbuff[14][28] ), 
        .D(\gbuff[15][28] ), .S0(n1447), .S1(n1426), .Y(n1365) );
  MX4X1 U526 ( .A(\gbuff[12][29] ), .B(\gbuff[13][29] ), .C(\gbuff[14][29] ), 
        .D(\gbuff[15][29] ), .S0(n1448), .S1(n1427), .Y(n1375) );
  MX4X1 U527 ( .A(\gbuff[12][30] ), .B(\gbuff[13][30] ), .C(\gbuff[14][30] ), 
        .D(\gbuff[15][30] ), .S0(n1430), .S1(n1428), .Y(n1385) );
  MX4X1 U528 ( .A(\gbuff[12][31] ), .B(\gbuff[13][31] ), .C(\gbuff[14][31] ), 
        .D(\gbuff[15][31] ), .S0(n1429), .S1(n1428), .Y(n1395) );
  MXI2X1 U529 ( .A(n36), .B(n37), .S0(n1401), .Y(N47) );
  MXI4X1 U530 ( .A(n31), .B(n29), .C(n30), .D(n28), .S0(n1403), .S1(n1409), 
        .Y(n37) );
  MXI4X1 U531 ( .A(n35), .B(n33), .C(n34), .D(n32), .S0(n1404), .S1(n1407), 
        .Y(n36) );
  MX4X1 U532 ( .A(\gbuff[28][0] ), .B(\gbuff[29][0] ), .C(\gbuff[30][0] ), .D(
        \gbuff[31][0] ), .S0(n1431), .S1(n1428), .Y(n28) );
  MXI2X1 U533 ( .A(n46), .B(n47), .S0(n1402), .Y(N46) );
  MXI4X1 U534 ( .A(n41), .B(n39), .C(n40), .D(n38), .S0(n1403), .S1(n1613), 
        .Y(n47) );
  MXI4X1 U535 ( .A(n45), .B(n43), .C(n44), .D(n42), .S0(n1404), .S1(n1408), 
        .Y(n46) );
  MX4X1 U536 ( .A(\gbuff[28][1] ), .B(\gbuff[29][1] ), .C(\gbuff[30][1] ), .D(
        \gbuff[31][1] ), .S0(n1431), .S1(n1427), .Y(n38) );
  MXI2X1 U537 ( .A(n56), .B(n57), .S0(N14), .Y(N45) );
  MXI4X1 U538 ( .A(n51), .B(n49), .C(n50), .D(n48), .S0(n1404), .S1(n1407), 
        .Y(n57) );
  MXI4X1 U539 ( .A(n55), .B(n53), .C(n54), .D(n52), .S0(n1404), .S1(n1407), 
        .Y(n56) );
  MX4X1 U540 ( .A(\gbuff[28][2] ), .B(\gbuff[29][2] ), .C(\gbuff[30][2] ), .D(
        \gbuff[31][2] ), .S0(n1432), .S1(n1411), .Y(n48) );
  MXI2X1 U541 ( .A(n66), .B(n67), .S0(N14), .Y(N44) );
  MXI4X1 U542 ( .A(n61), .B(n59), .C(n60), .D(n58), .S0(n1404), .S1(n1407), 
        .Y(n67) );
  MXI4X1 U543 ( .A(n65), .B(n63), .C(n64), .D(n62), .S0(n1404), .S1(n1407), 
        .Y(n66) );
  MX4X1 U544 ( .A(\gbuff[28][3] ), .B(\gbuff[29][3] ), .C(\gbuff[30][3] ), .D(
        \gbuff[31][3] ), .S0(n1433), .S1(n1412), .Y(n58) );
  MXI2X1 U545 ( .A(n76), .B(n77), .S0(N14), .Y(N43) );
  MXI4X1 U546 ( .A(n71), .B(n69), .C(n70), .D(n68), .S0(n1404), .S1(n1407), 
        .Y(n77) );
  MXI4X1 U547 ( .A(n75), .B(n73), .C(n74), .D(n72), .S0(n1404), .S1(n1407), 
        .Y(n76) );
  MX4X1 U548 ( .A(\gbuff[28][4] ), .B(\gbuff[29][4] ), .C(\gbuff[30][4] ), .D(
        \gbuff[31][4] ), .S0(n1433), .S1(n1412), .Y(n68) );
  MXI2X1 U549 ( .A(n86), .B(n87), .S0(N14), .Y(N42) );
  MXI4X1 U550 ( .A(n81), .B(n79), .C(n80), .D(n78), .S0(n1404), .S1(n1407), 
        .Y(n87) );
  MXI4X1 U551 ( .A(n85), .B(n83), .C(n84), .D(n82), .S0(n1404), .S1(n1407), 
        .Y(n86) );
  MX4X1 U552 ( .A(\gbuff[28][5] ), .B(\gbuff[29][5] ), .C(\gbuff[30][5] ), .D(
        \gbuff[31][5] ), .S0(n1434), .S1(n1424), .Y(n78) );
  MXI2X1 U553 ( .A(n96), .B(n97), .S0(N14), .Y(N41) );
  MXI4X1 U554 ( .A(n91), .B(n89), .C(n90), .D(n88), .S0(n1404), .S1(n1407), 
        .Y(n97) );
  MXI4X1 U555 ( .A(n95), .B(n93), .C(n94), .D(n92), .S0(n1404), .S1(n1407), 
        .Y(n96) );
  MX4X1 U556 ( .A(\gbuff[28][6] ), .B(\gbuff[29][6] ), .C(\gbuff[30][6] ), .D(
        \gbuff[31][6] ), .S0(n1435), .S1(n1413), .Y(n88) );
  MXI2X1 U557 ( .A(n112), .B(n114), .S0(N14), .Y(N40) );
  MXI4X1 U558 ( .A(n101), .B(n99), .C(n100), .D(n98), .S0(n1404), .S1(n1407), 
        .Y(n114) );
  MXI4X1 U559 ( .A(n110), .B(n106), .C(n108), .D(n104), .S0(n1404), .S1(n1407), 
        .Y(n112) );
  MX4X1 U560 ( .A(\gbuff[28][7] ), .B(\gbuff[29][7] ), .C(\gbuff[30][7] ), .D(
        \gbuff[31][7] ), .S0(n1435), .S1(n1413), .Y(n98) );
  MXI2X1 U561 ( .A(n127), .B(n1170), .S0(n1401), .Y(N39) );
  MXI4X1 U562 ( .A(n122), .B(n119), .C(n121), .D(n116), .S0(n1405), .S1(n1408), 
        .Y(n1170) );
  MXI4X1 U563 ( .A(n126), .B(n124), .C(n125), .D(n123), .S0(n1405), .S1(n1408), 
        .Y(n127) );
  MX4X1 U564 ( .A(\gbuff[28][8] ), .B(\gbuff[29][8] ), .C(\gbuff[30][8] ), .D(
        \gbuff[31][8] ), .S0(n1436), .S1(n1414), .Y(n116) );
  MXI2X1 U565 ( .A(n1179), .B(n1180), .S0(n1401), .Y(N38) );
  MXI4X1 U566 ( .A(n1174), .B(n1172), .C(n1173), .D(n1171), .S0(n1405), .S1(
        n1408), .Y(n1180) );
  MXI4X1 U567 ( .A(n1178), .B(n1176), .C(n1177), .D(n1175), .S0(n1405), .S1(
        n1408), .Y(n1179) );
  MX4X1 U568 ( .A(\gbuff[28][9] ), .B(\gbuff[29][9] ), .C(\gbuff[30][9] ), .D(
        \gbuff[31][9] ), .S0(n1436), .S1(n1414), .Y(n1171) );
  MXI2X1 U569 ( .A(n1189), .B(n1190), .S0(n1401), .Y(N37) );
  MXI4X1 U570 ( .A(n1184), .B(n1182), .C(n1183), .D(n1181), .S0(n1405), .S1(
        n1408), .Y(n1190) );
  MXI4X1 U571 ( .A(n1188), .B(n1186), .C(n1187), .D(n1185), .S0(n1405), .S1(
        n1408), .Y(n1189) );
  MX4X1 U572 ( .A(\gbuff[28][10] ), .B(\gbuff[29][10] ), .C(\gbuff[30][10] ), 
        .D(\gbuff[31][10] ), .S0(n1437), .S1(n1415), .Y(n1181) );
  MXI2X1 U573 ( .A(n1199), .B(n1200), .S0(n1401), .Y(N36) );
  MXI4X1 U574 ( .A(n1194), .B(n1192), .C(n1193), .D(n1191), .S0(n1405), .S1(
        n1408), .Y(n1200) );
  MXI4X1 U575 ( .A(n1198), .B(n1196), .C(n1197), .D(n1195), .S0(n1405), .S1(
        n1408), .Y(n1199) );
  MX4X1 U576 ( .A(\gbuff[28][11] ), .B(\gbuff[29][11] ), .C(\gbuff[30][11] ), 
        .D(\gbuff[31][11] ), .S0(n1438), .S1(n1416), .Y(n1191) );
  MXI2X1 U577 ( .A(n1209), .B(n1210), .S0(n1401), .Y(N35) );
  MXI4X1 U578 ( .A(n1204), .B(n1202), .C(n1203), .D(n1201), .S0(n1405), .S1(
        n1408), .Y(n1210) );
  MXI4X1 U579 ( .A(n1208), .B(n1206), .C(n1207), .D(n1205), .S0(n1405), .S1(
        n1408), .Y(n1209) );
  MX4X1 U580 ( .A(\gbuff[28][12] ), .B(\gbuff[29][12] ), .C(\gbuff[30][12] ), 
        .D(\gbuff[31][12] ), .S0(n1438), .S1(n1416), .Y(n1201) );
  MXI2X1 U581 ( .A(n1219), .B(n1220), .S0(n1401), .Y(N34) );
  MXI4X1 U582 ( .A(n1214), .B(n1212), .C(n1213), .D(n1211), .S0(n1405), .S1(
        n1408), .Y(n1220) );
  MXI4X1 U583 ( .A(n1218), .B(n1216), .C(n1217), .D(n1215), .S0(n1405), .S1(
        n1408), .Y(n1219) );
  MX4X1 U584 ( .A(\gbuff[28][13] ), .B(\gbuff[29][13] ), .C(\gbuff[30][13] ), 
        .D(\gbuff[31][13] ), .S0(n1439), .S1(n1417), .Y(n1211) );
  MXI2X1 U585 ( .A(n1229), .B(n1230), .S0(n1401), .Y(N33) );
  MXI4X1 U586 ( .A(n1224), .B(n1222), .C(n1223), .D(n1221), .S0(N13), .S1(
        n1409), .Y(n1230) );
  MXI4X1 U587 ( .A(n1228), .B(n1226), .C(n1227), .D(n1225), .S0(n1405), .S1(
        n1409), .Y(n1229) );
  MX4X1 U588 ( .A(\gbuff[28][14] ), .B(\gbuff[29][14] ), .C(\gbuff[30][14] ), 
        .D(\gbuff[31][14] ), .S0(n1439), .S1(n1417), .Y(n1221) );
  MXI2X1 U589 ( .A(n1239), .B(n1240), .S0(n1401), .Y(N32) );
  MXI4X1 U590 ( .A(n1234), .B(n1232), .C(n1233), .D(n1231), .S0(N13), .S1(
        n1409), .Y(n1240) );
  MXI4X1 U591 ( .A(n1238), .B(n1236), .C(n1237), .D(n1235), .S0(n1405), .S1(
        n1409), .Y(n1239) );
  MX4X1 U592 ( .A(\gbuff[28][15] ), .B(\gbuff[29][15] ), .C(\gbuff[30][15] ), 
        .D(\gbuff[31][15] ), .S0(n1440), .S1(n1418), .Y(n1231) );
  MXI2X1 U593 ( .A(n1249), .B(n1250), .S0(n1401), .Y(N31) );
  MXI4X1 U594 ( .A(n1244), .B(n1242), .C(n1243), .D(n1241), .S0(N13), .S1(
        n1409), .Y(n1250) );
  MXI4X1 U595 ( .A(n1248), .B(n1246), .C(n1247), .D(n1245), .S0(n1405), .S1(
        n1409), .Y(n1249) );
  MX4X1 U596 ( .A(\gbuff[28][16] ), .B(\gbuff[29][16] ), .C(\gbuff[30][16] ), 
        .D(\gbuff[31][16] ), .S0(n1441), .S1(n1419), .Y(n1241) );
  MXI2X1 U597 ( .A(n1259), .B(n1260), .S0(n1401), .Y(N30) );
  MXI4X1 U598 ( .A(n1254), .B(n1252), .C(n1253), .D(n1251), .S0(N13), .S1(
        n1409), .Y(n1260) );
  MXI4X1 U599 ( .A(n1258), .B(n1256), .C(n1257), .D(n1255), .S0(n1405), .S1(
        n1409), .Y(n1259) );
  MX4X1 U600 ( .A(\gbuff[28][17] ), .B(\gbuff[29][17] ), .C(\gbuff[30][17] ), 
        .D(\gbuff[31][17] ), .S0(n1441), .S1(n1419), .Y(n1251) );
  MXI2X1 U601 ( .A(n1269), .B(n1270), .S0(n1401), .Y(N29) );
  MXI4X1 U602 ( .A(n1264), .B(n1262), .C(n1263), .D(n1261), .S0(N13), .S1(
        n1409), .Y(n1270) );
  MXI4X1 U603 ( .A(n1268), .B(n1266), .C(n1267), .D(n1265), .S0(n1406), .S1(
        n1409), .Y(n1269) );
  MX4X1 U604 ( .A(\gbuff[28][18] ), .B(\gbuff[29][18] ), .C(\gbuff[30][18] ), 
        .D(\gbuff[31][18] ), .S0(n1442), .S1(n1420), .Y(n1261) );
  MXI2X1 U605 ( .A(n1279), .B(n1280), .S0(n1401), .Y(N28) );
  MXI4X1 U606 ( .A(n1274), .B(n1272), .C(n1273), .D(n1271), .S0(N13), .S1(
        n1409), .Y(n1280) );
  MXI4X1 U607 ( .A(n1278), .B(n1276), .C(n1277), .D(n1275), .S0(n1403), .S1(
        n1409), .Y(n1279) );
  MX4X1 U608 ( .A(\gbuff[28][19] ), .B(\gbuff[29][19] ), .C(\gbuff[30][19] ), 
        .D(\gbuff[31][19] ), .S0(n1443), .S1(n1421), .Y(n1271) );
  MXI2X1 U609 ( .A(n1289), .B(n1290), .S0(n1402), .Y(N27) );
  MXI4X1 U610 ( .A(n1284), .B(n1282), .C(n1283), .D(n1281), .S0(n1406), .S1(
        n1408), .Y(n1290) );
  MXI4X1 U611 ( .A(n1288), .B(n1286), .C(n1287), .D(n1285), .S0(n1406), .S1(
        n1408), .Y(n1289) );
  MX4X1 U612 ( .A(\gbuff[28][20] ), .B(\gbuff[29][20] ), .C(\gbuff[30][20] ), 
        .D(\gbuff[31][20] ), .S0(n1443), .S1(n1421), .Y(n1281) );
  MXI2X1 U613 ( .A(n1299), .B(n1300), .S0(n1402), .Y(N26) );
  MXI4X1 U614 ( .A(n1294), .B(n1292), .C(n1293), .D(n1291), .S0(n1406), .S1(
        n1409), .Y(n1300) );
  MXI4X1 U615 ( .A(n1298), .B(n1296), .C(n1297), .D(n1295), .S0(n1406), .S1(
        n1409), .Y(n1299) );
  MX4X1 U616 ( .A(\gbuff[28][21] ), .B(\gbuff[29][21] ), .C(\gbuff[30][21] ), 
        .D(\gbuff[31][21] ), .S0(n1444), .S1(n1422), .Y(n1291) );
  MXI2X1 U617 ( .A(n1309), .B(n1310), .S0(n1402), .Y(N25) );
  MXI4X1 U618 ( .A(n1304), .B(n1302), .C(n1303), .D(n1301), .S0(n1406), .S1(
        n1407), .Y(n1310) );
  MXI4X1 U619 ( .A(n1308), .B(n1306), .C(n1307), .D(n1305), .S0(n1406), .S1(
        n1407), .Y(n1309) );
  MX4X1 U620 ( .A(\gbuff[28][22] ), .B(\gbuff[29][22] ), .C(\gbuff[30][22] ), 
        .D(\gbuff[31][22] ), .S0(n1444), .S1(n1422), .Y(n1301) );
  MXI2X1 U621 ( .A(n1319), .B(n1320), .S0(n1402), .Y(N24) );
  MXI4X1 U622 ( .A(n1314), .B(n1312), .C(n1313), .D(n1311), .S0(n1406), .S1(
        n1408), .Y(n1320) );
  MXI4X1 U623 ( .A(n1318), .B(n1316), .C(n1317), .D(n1315), .S0(n1406), .S1(
        n1613), .Y(n1319) );
  MX4X1 U624 ( .A(\gbuff[28][23] ), .B(\gbuff[29][23] ), .C(\gbuff[30][23] ), 
        .D(\gbuff[31][23] ), .S0(n1445), .S1(n1423), .Y(n1311) );
  MXI2X1 U625 ( .A(n1329), .B(n1330), .S0(n1402), .Y(N23) );
  MXI4X1 U626 ( .A(n1324), .B(n1322), .C(n1323), .D(n1321), .S0(n1406), .S1(
        n1407), .Y(n1330) );
  MXI4X1 U627 ( .A(n1328), .B(n1326), .C(n1327), .D(n1325), .S0(n1406), .S1(
        n1408), .Y(n1329) );
  MX4X1 U628 ( .A(\gbuff[28][24] ), .B(\gbuff[29][24] ), .C(\gbuff[30][24] ), 
        .D(\gbuff[31][24] ), .S0(n1446), .S1(n1424), .Y(n1321) );
  MXI2X1 U629 ( .A(n1339), .B(n1340), .S0(n1402), .Y(N22) );
  MXI4X1 U630 ( .A(n1334), .B(n1332), .C(n1333), .D(n1331), .S0(n1406), .S1(
        n1408), .Y(n1340) );
  MXI4X1 U631 ( .A(n1338), .B(n1336), .C(n1337), .D(n1335), .S0(n1406), .S1(
        n1409), .Y(n1339) );
  MX4X1 U632 ( .A(\gbuff[28][25] ), .B(\gbuff[29][25] ), .C(\gbuff[30][25] ), 
        .D(\gbuff[31][25] ), .S0(n1446), .S1(n1424), .Y(n1331) );
  MXI2X1 U633 ( .A(n1349), .B(n1350), .S0(n1402), .Y(N21) );
  MXI4X1 U634 ( .A(n1344), .B(n1342), .C(n1343), .D(n1341), .S0(n1403), .S1(
        n1613), .Y(n1350) );
  MXI4X1 U635 ( .A(n1348), .B(n1346), .C(n1347), .D(n1345), .S0(n1403), .S1(
        n1407), .Y(n1349) );
  MX4X1 U636 ( .A(\gbuff[28][26] ), .B(\gbuff[29][26] ), .C(\gbuff[30][26] ), 
        .D(\gbuff[31][26] ), .S0(N10), .S1(n1425), .Y(n1341) );
  MXI2X1 U637 ( .A(n1359), .B(n1360), .S0(n1402), .Y(N20) );
  MXI4X1 U638 ( .A(n1354), .B(n1352), .C(n1353), .D(n1351), .S0(n1403), .S1(
        n1613), .Y(n1360) );
  MXI4X1 U639 ( .A(n1358), .B(n1356), .C(n1357), .D(n1355), .S0(n1404), .S1(
        n1613), .Y(n1359) );
  MX4X1 U640 ( .A(\gbuff[28][27] ), .B(\gbuff[29][27] ), .C(\gbuff[30][27] ), 
        .D(\gbuff[31][27] ), .S0(N10), .S1(n1425), .Y(n1351) );
  MXI2X1 U641 ( .A(n1369), .B(n1370), .S0(n1402), .Y(N19) );
  MXI4X1 U642 ( .A(n1364), .B(n1362), .C(n1363), .D(n1361), .S0(n1403), .S1(
        n1613), .Y(n1370) );
  MXI4X1 U643 ( .A(n1368), .B(n1366), .C(n1367), .D(n1365), .S0(n1404), .S1(
        n1409), .Y(n1369) );
  MX4X1 U644 ( .A(\gbuff[28][28] ), .B(\gbuff[29][28] ), .C(\gbuff[30][28] ), 
        .D(\gbuff[31][28] ), .S0(n1447), .S1(n1426), .Y(n1361) );
  MXI2X1 U645 ( .A(n1379), .B(n1380), .S0(n1402), .Y(N18) );
  MXI4X1 U646 ( .A(n1374), .B(n1372), .C(n1373), .D(n1371), .S0(n1403), .S1(
        n1613), .Y(n1380) );
  MXI4X1 U647 ( .A(n1378), .B(n1376), .C(n1377), .D(n1375), .S0(n1406), .S1(
        n1407), .Y(n1379) );
  MX4X1 U648 ( .A(\gbuff[28][29] ), .B(\gbuff[29][29] ), .C(\gbuff[30][29] ), 
        .D(\gbuff[31][29] ), .S0(n1448), .S1(n1427), .Y(n1371) );
  MXI2X1 U649 ( .A(n1389), .B(n1390), .S0(n1402), .Y(N17) );
  MXI4X1 U650 ( .A(n1384), .B(n1382), .C(n1383), .D(n1381), .S0(n1403), .S1(
        n1613), .Y(n1390) );
  MXI4X1 U651 ( .A(n1388), .B(n1386), .C(n1387), .D(n1385), .S0(N13), .S1(
        n1408), .Y(n1389) );
  MX4X1 U652 ( .A(\gbuff[28][30] ), .B(\gbuff[29][30] ), .C(\gbuff[30][30] ), 
        .D(\gbuff[31][30] ), .S0(n1448), .S1(n1427), .Y(n1381) );
  MXI2X1 U653 ( .A(n1399), .B(n1400), .S0(n1402), .Y(N16) );
  MXI4X1 U654 ( .A(n1394), .B(n1392), .C(n1393), .D(n1391), .S0(n1403), .S1(
        n1613), .Y(n1400) );
  MXI4X1 U655 ( .A(n1398), .B(n1396), .C(n1397), .D(n1395), .S0(N13), .S1(
        n1409), .Y(n1399) );
  MX4X1 U656 ( .A(\gbuff[28][31] ), .B(\gbuff[29][31] ), .C(\gbuff[30][31] ), 
        .D(\gbuff[31][31] ), .S0(n1430), .S1(n1428), .Y(n1391) );
  OAI2BB2XL U657 ( .B0(n1606), .B1(n1512), .A0N(\gbuff[0][0] ), .A1N(n1608), 
        .Y(n146) );
  OAI2BB2XL U658 ( .B0(n1607), .B1(n1510), .A0N(\gbuff[0][1] ), .A1N(n1606), 
        .Y(n147) );
  OAI2BB2XL U659 ( .B0(n1606), .B1(n1508), .A0N(\gbuff[0][2] ), .A1N(n1606), 
        .Y(n148) );
  OAI2BB2XL U660 ( .B0(n1606), .B1(n1506), .A0N(\gbuff[0][3] ), .A1N(n1608), 
        .Y(n149) );
  OAI2BB2XL U661 ( .B0(n1607), .B1(n1504), .A0N(\gbuff[0][4] ), .A1N(n1608), 
        .Y(n150) );
  OAI2BB2XL U662 ( .B0(n1606), .B1(n1502), .A0N(\gbuff[0][5] ), .A1N(n1608), 
        .Y(n151) );
  OAI2BB2XL U663 ( .B0(n1607), .B1(n1500), .A0N(\gbuff[0][6] ), .A1N(n1608), 
        .Y(n152) );
  OAI2BB2XL U664 ( .B0(n1606), .B1(n1498), .A0N(\gbuff[0][7] ), .A1N(n1608), 
        .Y(n153) );
  OAI2BB2XL U665 ( .B0(n1607), .B1(n1496), .A0N(\gbuff[0][8] ), .A1N(n1608), 
        .Y(n154) );
  OAI2BB2XL U666 ( .B0(n1606), .B1(n1494), .A0N(\gbuff[0][9] ), .A1N(n1608), 
        .Y(n155) );
  OAI2BB2XL U667 ( .B0(n1607), .B1(n1492), .A0N(\gbuff[0][10] ), .A1N(n1608), 
        .Y(n156) );
  OAI2BB2XL U668 ( .B0(n1606), .B1(n1490), .A0N(\gbuff[0][11] ), .A1N(n1608), 
        .Y(n157) );
  OAI2BB2XL U669 ( .B0(n1607), .B1(n1488), .A0N(\gbuff[0][12] ), .A1N(n1608), 
        .Y(n158) );
  OAI2BB2XL U670 ( .B0(n1606), .B1(n1486), .A0N(\gbuff[0][13] ), .A1N(n1608), 
        .Y(n159) );
  OAI2BB2XL U671 ( .B0(n1606), .B1(n1484), .A0N(\gbuff[0][14] ), .A1N(n1608), 
        .Y(n160) );
  OAI2BB2XL U672 ( .B0(n1606), .B1(n1482), .A0N(\gbuff[0][15] ), .A1N(n1607), 
        .Y(n161) );
  OAI2BB2XL U673 ( .B0(n1606), .B1(n1480), .A0N(\gbuff[0][16] ), .A1N(n1608), 
        .Y(n162) );
  OAI2BB2XL U674 ( .B0(n1606), .B1(n1478), .A0N(\gbuff[0][17] ), .A1N(n1607), 
        .Y(n163) );
  OAI2BB2XL U675 ( .B0(n1606), .B1(n1476), .A0N(\gbuff[0][18] ), .A1N(n1607), 
        .Y(n164) );
  OAI2BB2XL U676 ( .B0(n1606), .B1(n1474), .A0N(\gbuff[0][19] ), .A1N(n1607), 
        .Y(n165) );
  OAI2BB2XL U677 ( .B0(n1606), .B1(n1472), .A0N(\gbuff[0][20] ), .A1N(n1607), 
        .Y(n166) );
  OAI2BB2XL U678 ( .B0(n1606), .B1(n1470), .A0N(\gbuff[0][21] ), .A1N(n1607), 
        .Y(n167) );
  OAI2BB2XL U679 ( .B0(n1606), .B1(n1468), .A0N(\gbuff[0][22] ), .A1N(n1608), 
        .Y(n168) );
  OAI2BB2XL U680 ( .B0(n1607), .B1(n1466), .A0N(\gbuff[0][23] ), .A1N(n1607), 
        .Y(n169) );
  OAI2BB2XL U681 ( .B0(n1606), .B1(n1464), .A0N(\gbuff[0][24] ), .A1N(n1608), 
        .Y(n170) );
  OAI2BB2XL U682 ( .B0(n1607), .B1(n1462), .A0N(\gbuff[0][25] ), .A1N(n1608), 
        .Y(n171) );
  OAI2BB2XL U683 ( .B0(n1607), .B1(n1460), .A0N(\gbuff[0][26] ), .A1N(n1608), 
        .Y(n172) );
  OAI2BB2XL U684 ( .B0(n1607), .B1(n1458), .A0N(\gbuff[0][27] ), .A1N(n1608), 
        .Y(n173) );
  OAI2BB2XL U685 ( .B0(n1607), .B1(n1456), .A0N(\gbuff[0][28] ), .A1N(n1608), 
        .Y(n174) );
  OAI2BB2XL U686 ( .B0(n1607), .B1(n1454), .A0N(\gbuff[0][29] ), .A1N(n1608), 
        .Y(n175) );
  OAI2BB2XL U687 ( .B0(n1607), .B1(n1452), .A0N(\gbuff[0][30] ), .A1N(n1608), 
        .Y(n176) );
  OAI2BB2XL U688 ( .B0(n1607), .B1(n1450), .A0N(\gbuff[0][31] ), .A1N(n1606), 
        .Y(n177) );
  OAI2BB2XL U689 ( .B0(n1646), .B1(n1603), .A0N(\gbuff[1][0] ), .A1N(n1605), 
        .Y(n178) );
  OAI2BB2XL U690 ( .B0(n1645), .B1(n1603), .A0N(\gbuff[1][1] ), .A1N(n1605), 
        .Y(n179) );
  OAI2BB2XL U691 ( .B0(n1644), .B1(n1603), .A0N(\gbuff[1][2] ), .A1N(n1603), 
        .Y(n180) );
  OAI2BB2XL U692 ( .B0(n1643), .B1(n1603), .A0N(\gbuff[1][3] ), .A1N(n1605), 
        .Y(n181) );
  OAI2BB2XL U693 ( .B0(n1642), .B1(n1603), .A0N(\gbuff[1][4] ), .A1N(n1605), 
        .Y(n182) );
  OAI2BB2XL U694 ( .B0(n1641), .B1(n1603), .A0N(\gbuff[1][5] ), .A1N(n1605), 
        .Y(n183) );
  OAI2BB2XL U695 ( .B0(n1640), .B1(n1603), .A0N(\gbuff[1][6] ), .A1N(n1605), 
        .Y(n184) );
  OAI2BB2XL U696 ( .B0(n1639), .B1(n1603), .A0N(\gbuff[1][7] ), .A1N(n1605), 
        .Y(n185) );
  OAI2BB2XL U697 ( .B0(n1638), .B1(n1603), .A0N(\gbuff[1][8] ), .A1N(n1605), 
        .Y(n186) );
  OAI2BB2XL U698 ( .B0(n1637), .B1(n1603), .A0N(\gbuff[1][9] ), .A1N(n1605), 
        .Y(n187) );
  OAI2BB2XL U699 ( .B0(n1636), .B1(n1603), .A0N(\gbuff[1][10] ), .A1N(n1605), 
        .Y(n188) );
  OAI2BB2XL U700 ( .B0(n1635), .B1(n1603), .A0N(\gbuff[1][11] ), .A1N(n1605), 
        .Y(n189) );
  OAI2BB2XL U701 ( .B0(n1634), .B1(n1603), .A0N(\gbuff[1][12] ), .A1N(n1605), 
        .Y(n190) );
  OAI2BB2XL U702 ( .B0(n1633), .B1(n1603), .A0N(\gbuff[1][13] ), .A1N(n1605), 
        .Y(n191) );
  OAI2BB2XL U703 ( .B0(n1632), .B1(n1604), .A0N(\gbuff[1][14] ), .A1N(n1605), 
        .Y(n192) );
  OAI2BB2XL U704 ( .B0(n1631), .B1(n1603), .A0N(\gbuff[1][15] ), .A1N(n1604), 
        .Y(n193) );
  OAI2BB2XL U705 ( .B0(n1630), .B1(n1604), .A0N(\gbuff[1][16] ), .A1N(n1605), 
        .Y(n194) );
  OAI2BB2XL U706 ( .B0(n1629), .B1(n1603), .A0N(\gbuff[1][17] ), .A1N(n1604), 
        .Y(n195) );
  OAI2BB2XL U707 ( .B0(n1628), .B1(n1604), .A0N(\gbuff[1][18] ), .A1N(n1604), 
        .Y(n196) );
  OAI2BB2XL U708 ( .B0(n1627), .B1(n1603), .A0N(\gbuff[1][19] ), .A1N(n1604), 
        .Y(n197) );
  OAI2BB2XL U709 ( .B0(n1626), .B1(n1604), .A0N(\gbuff[1][20] ), .A1N(n1604), 
        .Y(n198) );
  OAI2BB2XL U710 ( .B0(n1625), .B1(n1603), .A0N(\gbuff[1][21] ), .A1N(n1604), 
        .Y(n199) );
  OAI2BB2XL U711 ( .B0(n1624), .B1(n1604), .A0N(\gbuff[1][22] ), .A1N(n1605), 
        .Y(n200) );
  OAI2BB2XL U712 ( .B0(n1623), .B1(n1604), .A0N(\gbuff[1][23] ), .A1N(n1604), 
        .Y(n201) );
  OAI2BB2XL U713 ( .B0(n1622), .B1(n1603), .A0N(\gbuff[1][24] ), .A1N(n1605), 
        .Y(n202) );
  OAI2BB2XL U714 ( .B0(n1621), .B1(n1604), .A0N(\gbuff[1][25] ), .A1N(n1605), 
        .Y(n203) );
  OAI2BB2XL U715 ( .B0(n1620), .B1(n1604), .A0N(\gbuff[1][26] ), .A1N(n1605), 
        .Y(n204) );
  OAI2BB2XL U716 ( .B0(n1619), .B1(n1604), .A0N(\gbuff[1][27] ), .A1N(n1605), 
        .Y(n205) );
  OAI2BB2XL U717 ( .B0(n1618), .B1(n1604), .A0N(\gbuff[1][28] ), .A1N(n1605), 
        .Y(n206) );
  OAI2BB2XL U718 ( .B0(n1617), .B1(n1604), .A0N(\gbuff[1][29] ), .A1N(n1605), 
        .Y(n207) );
  OAI2BB2XL U719 ( .B0(n1616), .B1(n1604), .A0N(\gbuff[1][30] ), .A1N(n1604), 
        .Y(n208) );
  OAI2BB2XL U720 ( .B0(n1615), .B1(n1604), .A0N(\gbuff[1][31] ), .A1N(n1603), 
        .Y(n209) );
  OAI2BB2XL U721 ( .B0(n1646), .B1(n1600), .A0N(\gbuff[2][0] ), .A1N(n1602), 
        .Y(n210) );
  OAI2BB2XL U722 ( .B0(n1645), .B1(n1600), .A0N(\gbuff[2][1] ), .A1N(n1602), 
        .Y(n211) );
  OAI2BB2XL U723 ( .B0(n1644), .B1(n1600), .A0N(\gbuff[2][2] ), .A1N(n1600), 
        .Y(n212) );
  OAI2BB2XL U724 ( .B0(n1643), .B1(n1600), .A0N(\gbuff[2][3] ), .A1N(n1602), 
        .Y(n213) );
  OAI2BB2XL U725 ( .B0(n1642), .B1(n1600), .A0N(\gbuff[2][4] ), .A1N(n1602), 
        .Y(n214) );
  OAI2BB2XL U726 ( .B0(n1641), .B1(n1600), .A0N(\gbuff[2][5] ), .A1N(n1602), 
        .Y(n215) );
  OAI2BB2XL U727 ( .B0(n1640), .B1(n1600), .A0N(\gbuff[2][6] ), .A1N(n1602), 
        .Y(n216) );
  OAI2BB2XL U728 ( .B0(n1639), .B1(n1600), .A0N(\gbuff[2][7] ), .A1N(n1602), 
        .Y(n217) );
  OAI2BB2XL U729 ( .B0(n1638), .B1(n1600), .A0N(\gbuff[2][8] ), .A1N(n1602), 
        .Y(n218) );
  OAI2BB2XL U730 ( .B0(n1637), .B1(n1600), .A0N(\gbuff[2][9] ), .A1N(n1602), 
        .Y(n219) );
  OAI2BB2XL U731 ( .B0(n1636), .B1(n1600), .A0N(\gbuff[2][10] ), .A1N(n1602), 
        .Y(n220) );
  OAI2BB2XL U732 ( .B0(n1635), .B1(n1600), .A0N(\gbuff[2][11] ), .A1N(n1602), 
        .Y(n221) );
  OAI2BB2XL U733 ( .B0(n1634), .B1(n1600), .A0N(\gbuff[2][12] ), .A1N(n1602), 
        .Y(n222) );
  OAI2BB2XL U734 ( .B0(n1633), .B1(n1600), .A0N(\gbuff[2][13] ), .A1N(n1602), 
        .Y(n223) );
  OAI2BB2XL U735 ( .B0(n1632), .B1(n1601), .A0N(\gbuff[2][14] ), .A1N(n1602), 
        .Y(n224) );
  OAI2BB2XL U736 ( .B0(n1631), .B1(n1600), .A0N(\gbuff[2][15] ), .A1N(n1601), 
        .Y(n225) );
  OAI2BB2XL U737 ( .B0(n1630), .B1(n1601), .A0N(\gbuff[2][16] ), .A1N(n1602), 
        .Y(n226) );
  OAI2BB2XL U738 ( .B0(n1629), .B1(n1600), .A0N(\gbuff[2][17] ), .A1N(n1601), 
        .Y(n227) );
  OAI2BB2XL U739 ( .B0(n1628), .B1(n1601), .A0N(\gbuff[2][18] ), .A1N(n1601), 
        .Y(n228) );
  OAI2BB2XL U740 ( .B0(n1627), .B1(n1600), .A0N(\gbuff[2][19] ), .A1N(n1601), 
        .Y(n229) );
  OAI2BB2XL U741 ( .B0(n1626), .B1(n1601), .A0N(\gbuff[2][20] ), .A1N(n1601), 
        .Y(n230) );
  OAI2BB2XL U742 ( .B0(n1625), .B1(n1600), .A0N(\gbuff[2][21] ), .A1N(n1601), 
        .Y(n231) );
  OAI2BB2XL U743 ( .B0(n1624), .B1(n1601), .A0N(\gbuff[2][22] ), .A1N(n1602), 
        .Y(n232) );
  OAI2BB2XL U744 ( .B0(n1623), .B1(n1601), .A0N(\gbuff[2][23] ), .A1N(n1601), 
        .Y(n233) );
  OAI2BB2XL U745 ( .B0(n1622), .B1(n1600), .A0N(\gbuff[2][24] ), .A1N(n1602), 
        .Y(n234) );
  OAI2BB2XL U746 ( .B0(n1621), .B1(n1601), .A0N(\gbuff[2][25] ), .A1N(n1602), 
        .Y(n235) );
  OAI2BB2XL U747 ( .B0(n1620), .B1(n1601), .A0N(\gbuff[2][26] ), .A1N(n1602), 
        .Y(n236) );
  OAI2BB2XL U748 ( .B0(n1619), .B1(n1601), .A0N(\gbuff[2][27] ), .A1N(n1602), 
        .Y(n237) );
  OAI2BB2XL U749 ( .B0(n1618), .B1(n1601), .A0N(\gbuff[2][28] ), .A1N(n1602), 
        .Y(n238) );
  OAI2BB2XL U750 ( .B0(n1617), .B1(n1601), .A0N(\gbuff[2][29] ), .A1N(n1602), 
        .Y(n239) );
  OAI2BB2XL U751 ( .B0(n1616), .B1(n1601), .A0N(\gbuff[2][30] ), .A1N(n1601), 
        .Y(n240) );
  OAI2BB2XL U752 ( .B0(n1615), .B1(n1601), .A0N(\gbuff[2][31] ), .A1N(n1600), 
        .Y(n241) );
  OAI2BB2XL U753 ( .B0(n1646), .B1(n1597), .A0N(\gbuff[3][0] ), .A1N(n1599), 
        .Y(n242) );
  OAI2BB2XL U754 ( .B0(n1645), .B1(n1597), .A0N(\gbuff[3][1] ), .A1N(n1599), 
        .Y(n243) );
  OAI2BB2XL U755 ( .B0(n1644), .B1(n1597), .A0N(\gbuff[3][2] ), .A1N(n1597), 
        .Y(n244) );
  OAI2BB2XL U756 ( .B0(n1643), .B1(n1597), .A0N(\gbuff[3][3] ), .A1N(n1599), 
        .Y(n245) );
  OAI2BB2XL U757 ( .B0(n1642), .B1(n1597), .A0N(\gbuff[3][4] ), .A1N(n1599), 
        .Y(n246) );
  OAI2BB2XL U758 ( .B0(n1641), .B1(n1597), .A0N(\gbuff[3][5] ), .A1N(n1599), 
        .Y(n247) );
  OAI2BB2XL U759 ( .B0(n1640), .B1(n1597), .A0N(\gbuff[3][6] ), .A1N(n1599), 
        .Y(n248) );
  OAI2BB2XL U760 ( .B0(n1639), .B1(n1597), .A0N(\gbuff[3][7] ), .A1N(n1599), 
        .Y(n249) );
  OAI2BB2XL U761 ( .B0(n1638), .B1(n1597), .A0N(\gbuff[3][8] ), .A1N(n1599), 
        .Y(n250) );
  OAI2BB2XL U762 ( .B0(n1637), .B1(n1597), .A0N(\gbuff[3][9] ), .A1N(n1599), 
        .Y(n251) );
  OAI2BB2XL U763 ( .B0(n1636), .B1(n1597), .A0N(\gbuff[3][10] ), .A1N(n1599), 
        .Y(n252) );
  OAI2BB2XL U764 ( .B0(n1635), .B1(n1597), .A0N(\gbuff[3][11] ), .A1N(n1599), 
        .Y(n253) );
  OAI2BB2XL U765 ( .B0(n1634), .B1(n1597), .A0N(\gbuff[3][12] ), .A1N(n1599), 
        .Y(n254) );
  OAI2BB2XL U766 ( .B0(n1633), .B1(n1597), .A0N(\gbuff[3][13] ), .A1N(n1599), 
        .Y(n255) );
  OAI2BB2XL U767 ( .B0(n1632), .B1(n1598), .A0N(\gbuff[3][14] ), .A1N(n1599), 
        .Y(n256) );
  OAI2BB2XL U768 ( .B0(n1631), .B1(n1597), .A0N(\gbuff[3][15] ), .A1N(n1598), 
        .Y(n257) );
  OAI2BB2XL U769 ( .B0(n1630), .B1(n1598), .A0N(\gbuff[3][16] ), .A1N(n1599), 
        .Y(n258) );
  OAI2BB2XL U770 ( .B0(n1629), .B1(n1597), .A0N(\gbuff[3][17] ), .A1N(n1598), 
        .Y(n259) );
  OAI2BB2XL U771 ( .B0(n1628), .B1(n1598), .A0N(\gbuff[3][18] ), .A1N(n1598), 
        .Y(n260) );
  OAI2BB2XL U772 ( .B0(n1627), .B1(n1597), .A0N(\gbuff[3][19] ), .A1N(n1598), 
        .Y(n261) );
  OAI2BB2XL U773 ( .B0(n1626), .B1(n1598), .A0N(\gbuff[3][20] ), .A1N(n1598), 
        .Y(n262) );
  OAI2BB2XL U774 ( .B0(n1625), .B1(n1597), .A0N(\gbuff[3][21] ), .A1N(n1598), 
        .Y(n263) );
  OAI2BB2XL U775 ( .B0(n1624), .B1(n1598), .A0N(\gbuff[3][22] ), .A1N(n1599), 
        .Y(n264) );
  OAI2BB2XL U776 ( .B0(n1623), .B1(n1598), .A0N(\gbuff[3][23] ), .A1N(n1598), 
        .Y(n265) );
  OAI2BB2XL U777 ( .B0(n1622), .B1(n1597), .A0N(\gbuff[3][24] ), .A1N(n1599), 
        .Y(n266) );
  OAI2BB2XL U778 ( .B0(n1621), .B1(n1598), .A0N(\gbuff[3][25] ), .A1N(n1599), 
        .Y(n267) );
  OAI2BB2XL U779 ( .B0(n1620), .B1(n1598), .A0N(\gbuff[3][26] ), .A1N(n1599), 
        .Y(n268) );
  OAI2BB2XL U780 ( .B0(n1619), .B1(n1598), .A0N(\gbuff[3][27] ), .A1N(n1599), 
        .Y(n269) );
  OAI2BB2XL U781 ( .B0(n1618), .B1(n1598), .A0N(\gbuff[3][28] ), .A1N(n1599), 
        .Y(n270) );
  OAI2BB2XL U782 ( .B0(n1617), .B1(n1598), .A0N(\gbuff[3][29] ), .A1N(n1599), 
        .Y(n271) );
  OAI2BB2XL U783 ( .B0(n1616), .B1(n1598), .A0N(\gbuff[3][30] ), .A1N(n1598), 
        .Y(n272) );
  OAI2BB2XL U784 ( .B0(n1615), .B1(n1598), .A0N(\gbuff[3][31] ), .A1N(n1597), 
        .Y(n273) );
  OAI2BB2XL U785 ( .B0(n1646), .B1(n1594), .A0N(\gbuff[4][0] ), .A1N(n1596), 
        .Y(n274) );
  OAI2BB2XL U786 ( .B0(n1645), .B1(n1594), .A0N(\gbuff[4][1] ), .A1N(n1594), 
        .Y(n275) );
  OAI2BB2XL U787 ( .B0(n1644), .B1(n1594), .A0N(\gbuff[4][2] ), .A1N(n1596), 
        .Y(n276) );
  OAI2BB2XL U788 ( .B0(n1643), .B1(n1594), .A0N(\gbuff[4][3] ), .A1N(n1596), 
        .Y(n277) );
  OAI2BB2XL U789 ( .B0(n1642), .B1(n1594), .A0N(\gbuff[4][4] ), .A1N(n1594), 
        .Y(n278) );
  OAI2BB2XL U790 ( .B0(n1641), .B1(n1594), .A0N(\gbuff[4][5] ), .A1N(n1596), 
        .Y(n279) );
  OAI2BB2XL U791 ( .B0(n1640), .B1(n1594), .A0N(\gbuff[4][6] ), .A1N(n1596), 
        .Y(n280) );
  OAI2BB2XL U792 ( .B0(n1639), .B1(n1594), .A0N(\gbuff[4][7] ), .A1N(n1596), 
        .Y(n281) );
  OAI2BB2XL U793 ( .B0(n1638), .B1(n1594), .A0N(\gbuff[4][8] ), .A1N(n1596), 
        .Y(n282) );
  OAI2BB2XL U794 ( .B0(n1637), .B1(n1594), .A0N(\gbuff[4][9] ), .A1N(n1596), 
        .Y(n283) );
  OAI2BB2XL U795 ( .B0(n1636), .B1(n1594), .A0N(\gbuff[4][10] ), .A1N(n1596), 
        .Y(n284) );
  OAI2BB2XL U796 ( .B0(n1635), .B1(n1594), .A0N(\gbuff[4][11] ), .A1N(n1596), 
        .Y(n285) );
  OAI2BB2XL U797 ( .B0(n1634), .B1(n1594), .A0N(\gbuff[4][12] ), .A1N(n1596), 
        .Y(n286) );
  OAI2BB2XL U798 ( .B0(n1633), .B1(n1595), .A0N(\gbuff[4][13] ), .A1N(n1596), 
        .Y(n287) );
  OAI2BB2XL U799 ( .B0(n1632), .B1(n1594), .A0N(\gbuff[4][14] ), .A1N(n1596), 
        .Y(n288) );
  OAI2BB2XL U800 ( .B0(n1631), .B1(n1595), .A0N(\gbuff[4][15] ), .A1N(n1595), 
        .Y(n289) );
  OAI2BB2XL U801 ( .B0(n1630), .B1(n1594), .A0N(\gbuff[4][16] ), .A1N(n1596), 
        .Y(n290) );
  OAI2BB2XL U802 ( .B0(n1629), .B1(n1595), .A0N(\gbuff[4][17] ), .A1N(n1595), 
        .Y(n291) );
  OAI2BB2XL U803 ( .B0(n1628), .B1(n1594), .A0N(\gbuff[4][18] ), .A1N(n1595), 
        .Y(n292) );
  OAI2BB2XL U804 ( .B0(n1627), .B1(n1595), .A0N(\gbuff[4][19] ), .A1N(n1595), 
        .Y(n293) );
  OAI2BB2XL U805 ( .B0(n1626), .B1(n1594), .A0N(\gbuff[4][20] ), .A1N(n1595), 
        .Y(n294) );
  OAI2BB2XL U806 ( .B0(n1625), .B1(n1595), .A0N(\gbuff[4][21] ), .A1N(n1595), 
        .Y(n295) );
  OAI2BB2XL U807 ( .B0(n1624), .B1(n1594), .A0N(\gbuff[4][22] ), .A1N(n1596), 
        .Y(n296) );
  OAI2BB2XL U808 ( .B0(n1623), .B1(n1595), .A0N(\gbuff[4][23] ), .A1N(n1595), 
        .Y(n297) );
  OAI2BB2XL U809 ( .B0(n1622), .B1(n1595), .A0N(\gbuff[4][24] ), .A1N(n1596), 
        .Y(n298) );
  OAI2BB2XL U810 ( .B0(n1621), .B1(n1595), .A0N(\gbuff[4][25] ), .A1N(n1596), 
        .Y(n299) );
  OAI2BB2XL U811 ( .B0(n1620), .B1(n1595), .A0N(\gbuff[4][26] ), .A1N(n1596), 
        .Y(n300) );
  OAI2BB2XL U812 ( .B0(n1619), .B1(n1595), .A0N(\gbuff[4][27] ), .A1N(n1596), 
        .Y(n301) );
  OAI2BB2XL U813 ( .B0(n1618), .B1(n1595), .A0N(\gbuff[4][28] ), .A1N(n1596), 
        .Y(n302) );
  OAI2BB2XL U814 ( .B0(n1617), .B1(n1595), .A0N(\gbuff[4][29] ), .A1N(n1596), 
        .Y(n303) );
  OAI2BB2XL U815 ( .B0(n1616), .B1(n1595), .A0N(\gbuff[4][30] ), .A1N(n1594), 
        .Y(n304) );
  OAI2BB2XL U816 ( .B0(n1615), .B1(n1595), .A0N(\gbuff[4][31] ), .A1N(n1596), 
        .Y(n305) );
  OAI2BB2XL U817 ( .B0(n1646), .B1(n1591), .A0N(\gbuff[5][0] ), .A1N(n1593), 
        .Y(n306) );
  OAI2BB2XL U818 ( .B0(n1645), .B1(n1591), .A0N(\gbuff[5][1] ), .A1N(n1593), 
        .Y(n307) );
  OAI2BB2XL U819 ( .B0(n1644), .B1(n1591), .A0N(\gbuff[5][2] ), .A1N(n1591), 
        .Y(n308) );
  OAI2BB2XL U820 ( .B0(n1643), .B1(n1591), .A0N(\gbuff[5][3] ), .A1N(n1593), 
        .Y(n309) );
  OAI2BB2XL U821 ( .B0(n1642), .B1(n1591), .A0N(\gbuff[5][4] ), .A1N(n1593), 
        .Y(n310) );
  OAI2BB2XL U822 ( .B0(n1641), .B1(n1591), .A0N(\gbuff[5][5] ), .A1N(n1593), 
        .Y(n311) );
  OAI2BB2XL U823 ( .B0(n1640), .B1(n1591), .A0N(\gbuff[5][6] ), .A1N(n1593), 
        .Y(n312) );
  OAI2BB2XL U824 ( .B0(n1639), .B1(n1591), .A0N(\gbuff[5][7] ), .A1N(n1593), 
        .Y(n313) );
  OAI2BB2XL U825 ( .B0(n1638), .B1(n1591), .A0N(\gbuff[5][8] ), .A1N(n1593), 
        .Y(n314) );
  OAI2BB2XL U826 ( .B0(n1637), .B1(n1591), .A0N(\gbuff[5][9] ), .A1N(n1593), 
        .Y(n315) );
  OAI2BB2XL U827 ( .B0(n1636), .B1(n1591), .A0N(\gbuff[5][10] ), .A1N(n1593), 
        .Y(n316) );
  OAI2BB2XL U828 ( .B0(n1635), .B1(n1591), .A0N(\gbuff[5][11] ), .A1N(n1593), 
        .Y(n317) );
  OAI2BB2XL U829 ( .B0(n1634), .B1(n1591), .A0N(\gbuff[5][12] ), .A1N(n1593), 
        .Y(n318) );
  OAI2BB2XL U830 ( .B0(n1633), .B1(n1591), .A0N(\gbuff[5][13] ), .A1N(n1593), 
        .Y(n319) );
  OAI2BB2XL U831 ( .B0(n1632), .B1(n1592), .A0N(\gbuff[5][14] ), .A1N(n1593), 
        .Y(n320) );
  OAI2BB2XL U832 ( .B0(n1631), .B1(n1591), .A0N(\gbuff[5][15] ), .A1N(n1592), 
        .Y(n321) );
  OAI2BB2XL U833 ( .B0(n1630), .B1(n1592), .A0N(\gbuff[5][16] ), .A1N(n1593), 
        .Y(n322) );
  OAI2BB2XL U834 ( .B0(n1629), .B1(n1591), .A0N(\gbuff[5][17] ), .A1N(n1592), 
        .Y(n323) );
  OAI2BB2XL U835 ( .B0(n1628), .B1(n1592), .A0N(\gbuff[5][18] ), .A1N(n1592), 
        .Y(n324) );
  OAI2BB2XL U836 ( .B0(n1627), .B1(n1591), .A0N(\gbuff[5][19] ), .A1N(n1592), 
        .Y(n325) );
  OAI2BB2XL U837 ( .B0(n1626), .B1(n1592), .A0N(\gbuff[5][20] ), .A1N(n1592), 
        .Y(n326) );
  OAI2BB2XL U838 ( .B0(n1625), .B1(n1591), .A0N(\gbuff[5][21] ), .A1N(n1592), 
        .Y(n327) );
  OAI2BB2XL U839 ( .B0(n1624), .B1(n1592), .A0N(\gbuff[5][22] ), .A1N(n1593), 
        .Y(n328) );
  OAI2BB2XL U840 ( .B0(n1623), .B1(n1592), .A0N(\gbuff[5][23] ), .A1N(n1592), 
        .Y(n329) );
  OAI2BB2XL U841 ( .B0(n1622), .B1(n6), .A0N(\gbuff[5][24] ), .A1N(n1593), .Y(
        n330) );
  OAI2BB2XL U842 ( .B0(n1621), .B1(n1592), .A0N(\gbuff[5][25] ), .A1N(n1593), 
        .Y(n331) );
  OAI2BB2XL U843 ( .B0(n1620), .B1(n1592), .A0N(\gbuff[5][26] ), .A1N(n1593), 
        .Y(n332) );
  OAI2BB2XL U844 ( .B0(n1619), .B1(n1592), .A0N(\gbuff[5][27] ), .A1N(n1593), 
        .Y(n333) );
  OAI2BB2XL U845 ( .B0(n1618), .B1(n1592), .A0N(\gbuff[5][28] ), .A1N(n1593), 
        .Y(n334) );
  OAI2BB2XL U846 ( .B0(n1617), .B1(n1592), .A0N(\gbuff[5][29] ), .A1N(n1593), 
        .Y(n335) );
  OAI2BB2XL U847 ( .B0(n1616), .B1(n1592), .A0N(\gbuff[5][30] ), .A1N(n6), .Y(
        n336) );
  OAI2BB2XL U848 ( .B0(n1615), .B1(n1592), .A0N(\gbuff[5][31] ), .A1N(n1591), 
        .Y(n337) );
  OAI2BB2XL U849 ( .B0(n1512), .B1(n1588), .A0N(\gbuff[6][0] ), .A1N(n1590), 
        .Y(n338) );
  OAI2BB2XL U850 ( .B0(n1510), .B1(n1588), .A0N(\gbuff[6][1] ), .A1N(n7), .Y(
        n339) );
  OAI2BB2XL U851 ( .B0(n1508), .B1(n1588), .A0N(\gbuff[6][2] ), .A1N(n1588), 
        .Y(n340) );
  OAI2BB2XL U852 ( .B0(n1506), .B1(n1588), .A0N(\gbuff[6][3] ), .A1N(n1590), 
        .Y(n341) );
  OAI2BB2XL U853 ( .B0(n1504), .B1(n1588), .A0N(\gbuff[6][4] ), .A1N(n1590), 
        .Y(n342) );
  OAI2BB2XL U854 ( .B0(n1502), .B1(n1588), .A0N(\gbuff[6][5] ), .A1N(n1590), 
        .Y(n343) );
  OAI2BB2XL U855 ( .B0(n1500), .B1(n1588), .A0N(\gbuff[6][6] ), .A1N(n1590), 
        .Y(n344) );
  OAI2BB2XL U856 ( .B0(n1498), .B1(n1588), .A0N(\gbuff[6][7] ), .A1N(n1590), 
        .Y(n345) );
  OAI2BB2XL U857 ( .B0(n1496), .B1(n1588), .A0N(\gbuff[6][8] ), .A1N(n1590), 
        .Y(n346) );
  OAI2BB2XL U858 ( .B0(n1494), .B1(n1588), .A0N(\gbuff[6][9] ), .A1N(n1590), 
        .Y(n347) );
  OAI2BB2XL U859 ( .B0(n1492), .B1(n1588), .A0N(\gbuff[6][10] ), .A1N(n1590), 
        .Y(n348) );
  OAI2BB2XL U860 ( .B0(n1490), .B1(n1588), .A0N(\gbuff[6][11] ), .A1N(n1590), 
        .Y(n349) );
  OAI2BB2XL U861 ( .B0(n1488), .B1(n1588), .A0N(\gbuff[6][12] ), .A1N(n1590), 
        .Y(n350) );
  OAI2BB2XL U862 ( .B0(n1486), .B1(n1588), .A0N(\gbuff[6][13] ), .A1N(n1590), 
        .Y(n351) );
  OAI2BB2XL U863 ( .B0(n1484), .B1(n1589), .A0N(\gbuff[6][14] ), .A1N(n1590), 
        .Y(n352) );
  OAI2BB2XL U864 ( .B0(n1482), .B1(n1588), .A0N(\gbuff[6][15] ), .A1N(n1589), 
        .Y(n353) );
  OAI2BB2XL U865 ( .B0(n1480), .B1(n1589), .A0N(\gbuff[6][16] ), .A1N(n1590), 
        .Y(n354) );
  OAI2BB2XL U866 ( .B0(n1478), .B1(n1588), .A0N(\gbuff[6][17] ), .A1N(n1589), 
        .Y(n355) );
  OAI2BB2XL U867 ( .B0(n1476), .B1(n1589), .A0N(\gbuff[6][18] ), .A1N(n1589), 
        .Y(n356) );
  OAI2BB2XL U868 ( .B0(n1474), .B1(n1588), .A0N(\gbuff[6][19] ), .A1N(n1589), 
        .Y(n357) );
  OAI2BB2XL U869 ( .B0(n1472), .B1(n1589), .A0N(\gbuff[6][20] ), .A1N(n1589), 
        .Y(n358) );
  OAI2BB2XL U870 ( .B0(n1470), .B1(n1588), .A0N(\gbuff[6][21] ), .A1N(n1589), 
        .Y(n359) );
  OAI2BB2XL U871 ( .B0(n1468), .B1(n1589), .A0N(\gbuff[6][22] ), .A1N(n1590), 
        .Y(n360) );
  OAI2BB2XL U872 ( .B0(n1466), .B1(n1589), .A0N(\gbuff[6][23] ), .A1N(n1589), 
        .Y(n361) );
  OAI2BB2XL U873 ( .B0(n1464), .B1(n7), .A0N(\gbuff[6][24] ), .A1N(n1590), .Y(
        n362) );
  OAI2BB2XL U874 ( .B0(n1462), .B1(n1589), .A0N(\gbuff[6][25] ), .A1N(n1590), 
        .Y(n363) );
  OAI2BB2XL U875 ( .B0(n1460), .B1(n1589), .A0N(\gbuff[6][26] ), .A1N(n1590), 
        .Y(n364) );
  OAI2BB2XL U876 ( .B0(n1458), .B1(n1589), .A0N(\gbuff[6][27] ), .A1N(n1590), 
        .Y(n365) );
  OAI2BB2XL U877 ( .B0(n1456), .B1(n1589), .A0N(\gbuff[6][28] ), .A1N(n1590), 
        .Y(n366) );
  OAI2BB2XL U878 ( .B0(n1454), .B1(n1589), .A0N(\gbuff[6][29] ), .A1N(n1590), 
        .Y(n367) );
  OAI2BB2XL U879 ( .B0(n1452), .B1(n1589), .A0N(\gbuff[6][30] ), .A1N(n1590), 
        .Y(n368) );
  OAI2BB2XL U880 ( .B0(n1450), .B1(n1589), .A0N(\gbuff[6][31] ), .A1N(n1588), 
        .Y(n369) );
  OAI2BB2XL U881 ( .B0(n1511), .B1(n1585), .A0N(\gbuff[7][0] ), .A1N(n1587), 
        .Y(n370) );
  OAI2BB2XL U882 ( .B0(n1509), .B1(n1585), .A0N(\gbuff[7][1] ), .A1N(n8), .Y(
        n371) );
  OAI2BB2XL U883 ( .B0(n1507), .B1(n1585), .A0N(\gbuff[7][2] ), .A1N(n1585), 
        .Y(n372) );
  OAI2BB2XL U884 ( .B0(n1505), .B1(n1585), .A0N(\gbuff[7][3] ), .A1N(n1587), 
        .Y(n373) );
  OAI2BB2XL U885 ( .B0(n1503), .B1(n1585), .A0N(\gbuff[7][4] ), .A1N(n1587), 
        .Y(n374) );
  OAI2BB2XL U886 ( .B0(n1501), .B1(n1585), .A0N(\gbuff[7][5] ), .A1N(n1587), 
        .Y(n375) );
  OAI2BB2XL U887 ( .B0(n1499), .B1(n1585), .A0N(\gbuff[7][6] ), .A1N(n1587), 
        .Y(n376) );
  OAI2BB2XL U888 ( .B0(n1497), .B1(n1585), .A0N(\gbuff[7][7] ), .A1N(n1587), 
        .Y(n377) );
  OAI2BB2XL U889 ( .B0(n1495), .B1(n1585), .A0N(\gbuff[7][8] ), .A1N(n1587), 
        .Y(n378) );
  OAI2BB2XL U890 ( .B0(n1493), .B1(n1585), .A0N(\gbuff[7][9] ), .A1N(n1587), 
        .Y(n379) );
  OAI2BB2XL U891 ( .B0(n1491), .B1(n1585), .A0N(\gbuff[7][10] ), .A1N(n1587), 
        .Y(n380) );
  OAI2BB2XL U892 ( .B0(n1489), .B1(n1585), .A0N(\gbuff[7][11] ), .A1N(n1587), 
        .Y(n381) );
  OAI2BB2XL U893 ( .B0(n1487), .B1(n1585), .A0N(\gbuff[7][12] ), .A1N(n1587), 
        .Y(n382) );
  OAI2BB2XL U894 ( .B0(n1485), .B1(n1585), .A0N(\gbuff[7][13] ), .A1N(n1587), 
        .Y(n383) );
  OAI2BB2XL U895 ( .B0(n1483), .B1(n1586), .A0N(\gbuff[7][14] ), .A1N(n1587), 
        .Y(n384) );
  OAI2BB2XL U896 ( .B0(n1481), .B1(n1585), .A0N(\gbuff[7][15] ), .A1N(n1586), 
        .Y(n385) );
  OAI2BB2XL U897 ( .B0(n1479), .B1(n1586), .A0N(\gbuff[7][16] ), .A1N(n1587), 
        .Y(n386) );
  OAI2BB2XL U898 ( .B0(n1477), .B1(n1585), .A0N(\gbuff[7][17] ), .A1N(n1586), 
        .Y(n387) );
  OAI2BB2XL U899 ( .B0(n1475), .B1(n1586), .A0N(\gbuff[7][18] ), .A1N(n1586), 
        .Y(n388) );
  OAI2BB2XL U900 ( .B0(n1473), .B1(n1585), .A0N(\gbuff[7][19] ), .A1N(n1586), 
        .Y(n389) );
  OAI2BB2XL U901 ( .B0(n1471), .B1(n1586), .A0N(\gbuff[7][20] ), .A1N(n1586), 
        .Y(n390) );
  OAI2BB2XL U902 ( .B0(n1469), .B1(n1585), .A0N(\gbuff[7][21] ), .A1N(n1586), 
        .Y(n391) );
  OAI2BB2XL U903 ( .B0(n1467), .B1(n1586), .A0N(\gbuff[7][22] ), .A1N(n1587), 
        .Y(n392) );
  OAI2BB2XL U904 ( .B0(n1465), .B1(n1586), .A0N(\gbuff[7][23] ), .A1N(n1586), 
        .Y(n393) );
  OAI2BB2XL U905 ( .B0(n1463), .B1(n8), .A0N(\gbuff[7][24] ), .A1N(n1587), .Y(
        n394) );
  OAI2BB2XL U906 ( .B0(n1461), .B1(n1586), .A0N(\gbuff[7][25] ), .A1N(n1587), 
        .Y(n395) );
  OAI2BB2XL U907 ( .B0(n1459), .B1(n1586), .A0N(\gbuff[7][26] ), .A1N(n1587), 
        .Y(n396) );
  OAI2BB2XL U908 ( .B0(n1457), .B1(n1586), .A0N(\gbuff[7][27] ), .A1N(n1587), 
        .Y(n397) );
  OAI2BB2XL U909 ( .B0(n1455), .B1(n1586), .A0N(\gbuff[7][28] ), .A1N(n1587), 
        .Y(n398) );
  OAI2BB2XL U910 ( .B0(n1453), .B1(n1586), .A0N(\gbuff[7][29] ), .A1N(n1587), 
        .Y(n399) );
  OAI2BB2XL U911 ( .B0(n1451), .B1(n1586), .A0N(\gbuff[7][30] ), .A1N(n1587), 
        .Y(n400) );
  OAI2BB2XL U912 ( .B0(n1449), .B1(n1586), .A0N(\gbuff[7][31] ), .A1N(n1585), 
        .Y(n401) );
  OAI2BB2XL U913 ( .B0(n1512), .B1(n1582), .A0N(\gbuff[8][0] ), .A1N(n1584), 
        .Y(n402) );
  OAI2BB2XL U914 ( .B0(n1510), .B1(n1582), .A0N(\gbuff[8][1] ), .A1N(n1583), 
        .Y(n403) );
  OAI2BB2XL U915 ( .B0(n1508), .B1(n1582), .A0N(\gbuff[8][2] ), .A1N(n1582), 
        .Y(n404) );
  OAI2BB2XL U916 ( .B0(n1506), .B1(n1582), .A0N(\gbuff[8][3] ), .A1N(n1584), 
        .Y(n405) );
  OAI2BB2XL U917 ( .B0(n1504), .B1(n1582), .A0N(\gbuff[8][4] ), .A1N(n1584), 
        .Y(n406) );
  OAI2BB2XL U918 ( .B0(n1502), .B1(n1582), .A0N(\gbuff[8][5] ), .A1N(n1584), 
        .Y(n407) );
  OAI2BB2XL U919 ( .B0(n1500), .B1(n1582), .A0N(\gbuff[8][6] ), .A1N(n1584), 
        .Y(n408) );
  OAI2BB2XL U920 ( .B0(n1498), .B1(n1582), .A0N(\gbuff[8][7] ), .A1N(n1584), 
        .Y(n409) );
  OAI2BB2XL U921 ( .B0(n1496), .B1(n1582), .A0N(\gbuff[8][8] ), .A1N(n1584), 
        .Y(n410) );
  OAI2BB2XL U922 ( .B0(n1494), .B1(n1582), .A0N(\gbuff[8][9] ), .A1N(n1584), 
        .Y(n411) );
  OAI2BB2XL U923 ( .B0(n1492), .B1(n1582), .A0N(\gbuff[8][10] ), .A1N(n1584), 
        .Y(n412) );
  OAI2BB2XL U924 ( .B0(n1490), .B1(n1582), .A0N(\gbuff[8][11] ), .A1N(n1584), 
        .Y(n413) );
  OAI2BB2XL U925 ( .B0(n1488), .B1(n1582), .A0N(\gbuff[8][12] ), .A1N(n1584), 
        .Y(n414) );
  OAI2BB2XL U926 ( .B0(n1486), .B1(n1582), .A0N(\gbuff[8][13] ), .A1N(n1584), 
        .Y(n415) );
  OAI2BB2XL U927 ( .B0(n1484), .B1(n1583), .A0N(\gbuff[8][14] ), .A1N(n1584), 
        .Y(n416) );
  OAI2BB2XL U928 ( .B0(n1482), .B1(n1582), .A0N(\gbuff[8][15] ), .A1N(n1583), 
        .Y(n417) );
  OAI2BB2XL U929 ( .B0(n1480), .B1(n1583), .A0N(\gbuff[8][16] ), .A1N(n1584), 
        .Y(n418) );
  OAI2BB2XL U930 ( .B0(n1478), .B1(n1582), .A0N(\gbuff[8][17] ), .A1N(n1583), 
        .Y(n419) );
  OAI2BB2XL U931 ( .B0(n1476), .B1(n1583), .A0N(\gbuff[8][18] ), .A1N(n1583), 
        .Y(n420) );
  OAI2BB2XL U932 ( .B0(n1474), .B1(n1582), .A0N(\gbuff[8][19] ), .A1N(n1583), 
        .Y(n421) );
  OAI2BB2XL U933 ( .B0(n1472), .B1(n1583), .A0N(\gbuff[8][20] ), .A1N(n1583), 
        .Y(n422) );
  OAI2BB2XL U934 ( .B0(n1470), .B1(n1582), .A0N(\gbuff[8][21] ), .A1N(n1583), 
        .Y(n423) );
  OAI2BB2XL U935 ( .B0(n1468), .B1(n1583), .A0N(\gbuff[8][22] ), .A1N(n1584), 
        .Y(n424) );
  OAI2BB2XL U936 ( .B0(n1466), .B1(n1583), .A0N(\gbuff[8][23] ), .A1N(n1583), 
        .Y(n425) );
  OAI2BB2XL U937 ( .B0(n1464), .B1(n1582), .A0N(\gbuff[8][24] ), .A1N(n1584), 
        .Y(n426) );
  OAI2BB2XL U938 ( .B0(n1462), .B1(n1583), .A0N(\gbuff[8][25] ), .A1N(n1584), 
        .Y(n427) );
  OAI2BB2XL U939 ( .B0(n1460), .B1(n1583), .A0N(\gbuff[8][26] ), .A1N(n1584), 
        .Y(n428) );
  OAI2BB2XL U940 ( .B0(n1458), .B1(n1583), .A0N(\gbuff[8][27] ), .A1N(n1584), 
        .Y(n429) );
  OAI2BB2XL U941 ( .B0(n1456), .B1(n1583), .A0N(\gbuff[8][28] ), .A1N(n1584), 
        .Y(n430) );
  OAI2BB2XL U942 ( .B0(n1454), .B1(n1583), .A0N(\gbuff[8][29] ), .A1N(n1584), 
        .Y(n431) );
  OAI2BB2XL U943 ( .B0(n1452), .B1(n1583), .A0N(\gbuff[8][30] ), .A1N(n1584), 
        .Y(n432) );
  OAI2BB2XL U944 ( .B0(n1450), .B1(n1583), .A0N(\gbuff[8][31] ), .A1N(n1582), 
        .Y(n433) );
  OAI2BB2XL U945 ( .B0(n1512), .B1(n1579), .A0N(\gbuff[9][0] ), .A1N(n1581), 
        .Y(n434) );
  OAI2BB2XL U946 ( .B0(n1510), .B1(n1579), .A0N(\gbuff[9][1] ), .A1N(n1580), 
        .Y(n435) );
  OAI2BB2XL U947 ( .B0(n1508), .B1(n1579), .A0N(\gbuff[9][2] ), .A1N(n1579), 
        .Y(n436) );
  OAI2BB2XL U948 ( .B0(n1506), .B1(n1579), .A0N(\gbuff[9][3] ), .A1N(n1581), 
        .Y(n437) );
  OAI2BB2XL U949 ( .B0(n1504), .B1(n1579), .A0N(\gbuff[9][4] ), .A1N(n1581), 
        .Y(n438) );
  OAI2BB2XL U950 ( .B0(n1502), .B1(n1579), .A0N(\gbuff[9][5] ), .A1N(n1581), 
        .Y(n439) );
  OAI2BB2XL U951 ( .B0(n1500), .B1(n1579), .A0N(\gbuff[9][6] ), .A1N(n1581), 
        .Y(n440) );
  OAI2BB2XL U952 ( .B0(n1498), .B1(n1579), .A0N(\gbuff[9][7] ), .A1N(n1581), 
        .Y(n441) );
  OAI2BB2XL U953 ( .B0(n1496), .B1(n1579), .A0N(\gbuff[9][8] ), .A1N(n1581), 
        .Y(n442) );
  OAI2BB2XL U954 ( .B0(n1494), .B1(n1579), .A0N(\gbuff[9][9] ), .A1N(n1581), 
        .Y(n443) );
  OAI2BB2XL U955 ( .B0(n1492), .B1(n1579), .A0N(\gbuff[9][10] ), .A1N(n1581), 
        .Y(n444) );
  OAI2BB2XL U956 ( .B0(n1490), .B1(n1579), .A0N(\gbuff[9][11] ), .A1N(n1581), 
        .Y(n445) );
  OAI2BB2XL U957 ( .B0(n1488), .B1(n1579), .A0N(\gbuff[9][12] ), .A1N(n1581), 
        .Y(n446) );
  OAI2BB2XL U958 ( .B0(n1486), .B1(n1579), .A0N(\gbuff[9][13] ), .A1N(n1581), 
        .Y(n447) );
  OAI2BB2XL U959 ( .B0(n1484), .B1(n1580), .A0N(\gbuff[9][14] ), .A1N(n1581), 
        .Y(n448) );
  OAI2BB2XL U960 ( .B0(n1482), .B1(n1579), .A0N(\gbuff[9][15] ), .A1N(n1580), 
        .Y(n449) );
  OAI2BB2XL U961 ( .B0(n1480), .B1(n1580), .A0N(\gbuff[9][16] ), .A1N(n1581), 
        .Y(n450) );
  OAI2BB2XL U962 ( .B0(n1478), .B1(n1579), .A0N(\gbuff[9][17] ), .A1N(n1580), 
        .Y(n451) );
  OAI2BB2XL U963 ( .B0(n1476), .B1(n1580), .A0N(\gbuff[9][18] ), .A1N(n1580), 
        .Y(n452) );
  OAI2BB2XL U964 ( .B0(n1474), .B1(n1579), .A0N(\gbuff[9][19] ), .A1N(n1580), 
        .Y(n453) );
  OAI2BB2XL U965 ( .B0(n1472), .B1(n1580), .A0N(\gbuff[9][20] ), .A1N(n1580), 
        .Y(n454) );
  OAI2BB2XL U966 ( .B0(n1470), .B1(n1579), .A0N(\gbuff[9][21] ), .A1N(n1580), 
        .Y(n455) );
  OAI2BB2XL U967 ( .B0(n1468), .B1(n1580), .A0N(\gbuff[9][22] ), .A1N(n1581), 
        .Y(n456) );
  OAI2BB2XL U968 ( .B0(n1466), .B1(n1580), .A0N(\gbuff[9][23] ), .A1N(n1580), 
        .Y(n457) );
  OAI2BB2XL U969 ( .B0(n1464), .B1(n1579), .A0N(\gbuff[9][24] ), .A1N(n1581), 
        .Y(n458) );
  OAI2BB2XL U970 ( .B0(n1462), .B1(n1580), .A0N(\gbuff[9][25] ), .A1N(n1581), 
        .Y(n459) );
  OAI2BB2XL U971 ( .B0(n1460), .B1(n1580), .A0N(\gbuff[9][26] ), .A1N(n1581), 
        .Y(n460) );
  OAI2BB2XL U972 ( .B0(n1458), .B1(n1580), .A0N(\gbuff[9][27] ), .A1N(n1581), 
        .Y(n461) );
  OAI2BB2XL U973 ( .B0(n1456), .B1(n1580), .A0N(\gbuff[9][28] ), .A1N(n1581), 
        .Y(n462) );
  OAI2BB2XL U974 ( .B0(n1454), .B1(n1580), .A0N(\gbuff[9][29] ), .A1N(n1581), 
        .Y(n463) );
  OAI2BB2XL U975 ( .B0(n1452), .B1(n1580), .A0N(\gbuff[9][30] ), .A1N(n1581), 
        .Y(n464) );
  OAI2BB2XL U976 ( .B0(n1450), .B1(n1580), .A0N(\gbuff[9][31] ), .A1N(n1579), 
        .Y(n465) );
  OAI2BB2XL U977 ( .B0(n1512), .B1(n1576), .A0N(\gbuff[10][0] ), .A1N(n1578), 
        .Y(n466) );
  OAI2BB2XL U978 ( .B0(n1510), .B1(n1576), .A0N(\gbuff[10][1] ), .A1N(n1577), 
        .Y(n467) );
  OAI2BB2XL U979 ( .B0(n1508), .B1(n1576), .A0N(\gbuff[10][2] ), .A1N(n1576), 
        .Y(n468) );
  OAI2BB2XL U980 ( .B0(n1506), .B1(n1576), .A0N(\gbuff[10][3] ), .A1N(n1578), 
        .Y(n469) );
  OAI2BB2XL U981 ( .B0(n1504), .B1(n1576), .A0N(\gbuff[10][4] ), .A1N(n1578), 
        .Y(n470) );
  OAI2BB2XL U982 ( .B0(n1502), .B1(n1576), .A0N(\gbuff[10][5] ), .A1N(n1578), 
        .Y(n471) );
  OAI2BB2XL U983 ( .B0(n1500), .B1(n1576), .A0N(\gbuff[10][6] ), .A1N(n1578), 
        .Y(n472) );
  OAI2BB2XL U984 ( .B0(n1498), .B1(n1576), .A0N(\gbuff[10][7] ), .A1N(n1578), 
        .Y(n473) );
  OAI2BB2XL U985 ( .B0(n1496), .B1(n1576), .A0N(\gbuff[10][8] ), .A1N(n1578), 
        .Y(n474) );
  OAI2BB2XL U986 ( .B0(n1494), .B1(n1576), .A0N(\gbuff[10][9] ), .A1N(n1578), 
        .Y(n475) );
  OAI2BB2XL U987 ( .B0(n1492), .B1(n1576), .A0N(\gbuff[10][10] ), .A1N(n1578), 
        .Y(n476) );
  OAI2BB2XL U988 ( .B0(n1490), .B1(n1576), .A0N(\gbuff[10][11] ), .A1N(n1578), 
        .Y(n477) );
  OAI2BB2XL U989 ( .B0(n1488), .B1(n1576), .A0N(\gbuff[10][12] ), .A1N(n1578), 
        .Y(n478) );
  OAI2BB2XL U990 ( .B0(n1486), .B1(n1576), .A0N(\gbuff[10][13] ), .A1N(n1578), 
        .Y(n479) );
  OAI2BB2XL U991 ( .B0(n1484), .B1(n1577), .A0N(\gbuff[10][14] ), .A1N(n1578), 
        .Y(n480) );
  OAI2BB2XL U992 ( .B0(n1482), .B1(n1576), .A0N(\gbuff[10][15] ), .A1N(n1577), 
        .Y(n481) );
  OAI2BB2XL U993 ( .B0(n1480), .B1(n1577), .A0N(\gbuff[10][16] ), .A1N(n1578), 
        .Y(n482) );
  OAI2BB2XL U994 ( .B0(n1478), .B1(n1576), .A0N(\gbuff[10][17] ), .A1N(n1577), 
        .Y(n483) );
  OAI2BB2XL U995 ( .B0(n1476), .B1(n1577), .A0N(\gbuff[10][18] ), .A1N(n1577), 
        .Y(n484) );
  OAI2BB2XL U996 ( .B0(n1474), .B1(n1576), .A0N(\gbuff[10][19] ), .A1N(n1577), 
        .Y(n485) );
  OAI2BB2XL U997 ( .B0(n1472), .B1(n1577), .A0N(\gbuff[10][20] ), .A1N(n1577), 
        .Y(n486) );
  OAI2BB2XL U998 ( .B0(n1470), .B1(n1576), .A0N(\gbuff[10][21] ), .A1N(n1577), 
        .Y(n487) );
  OAI2BB2XL U999 ( .B0(n1468), .B1(n1577), .A0N(\gbuff[10][22] ), .A1N(n1578), 
        .Y(n488) );
  OAI2BB2XL U1000 ( .B0(n1466), .B1(n1577), .A0N(\gbuff[10][23] ), .A1N(n1577), 
        .Y(n489) );
  OAI2BB2XL U1001 ( .B0(n1464), .B1(n1576), .A0N(\gbuff[10][24] ), .A1N(n1578), 
        .Y(n490) );
  OAI2BB2XL U1002 ( .B0(n1462), .B1(n1577), .A0N(\gbuff[10][25] ), .A1N(n1578), 
        .Y(n491) );
  OAI2BB2XL U1003 ( .B0(n1460), .B1(n1577), .A0N(\gbuff[10][26] ), .A1N(n1578), 
        .Y(n492) );
  OAI2BB2XL U1004 ( .B0(n1458), .B1(n1577), .A0N(\gbuff[10][27] ), .A1N(n1578), 
        .Y(n493) );
  OAI2BB2XL U1005 ( .B0(n1456), .B1(n1577), .A0N(\gbuff[10][28] ), .A1N(n1578), 
        .Y(n494) );
  OAI2BB2XL U1006 ( .B0(n1454), .B1(n1577), .A0N(\gbuff[10][29] ), .A1N(n1578), 
        .Y(n495) );
  OAI2BB2XL U1007 ( .B0(n1452), .B1(n1577), .A0N(\gbuff[10][30] ), .A1N(n1578), 
        .Y(n496) );
  OAI2BB2XL U1008 ( .B0(n1450), .B1(n1577), .A0N(\gbuff[10][31] ), .A1N(n1576), 
        .Y(n497) );
  OAI2BB2XL U1009 ( .B0(n1512), .B1(n1573), .A0N(\gbuff[11][0] ), .A1N(n1575), 
        .Y(n498) );
  OAI2BB2XL U1010 ( .B0(n1510), .B1(n1573), .A0N(\gbuff[11][1] ), .A1N(n1574), 
        .Y(n499) );
  OAI2BB2XL U1011 ( .B0(n1508), .B1(n1573), .A0N(\gbuff[11][2] ), .A1N(n1573), 
        .Y(n500) );
  OAI2BB2XL U1012 ( .B0(n1506), .B1(n1573), .A0N(\gbuff[11][3] ), .A1N(n1575), 
        .Y(n501) );
  OAI2BB2XL U1013 ( .B0(n1504), .B1(n1573), .A0N(\gbuff[11][4] ), .A1N(n1575), 
        .Y(n502) );
  OAI2BB2XL U1014 ( .B0(n1502), .B1(n1573), .A0N(\gbuff[11][5] ), .A1N(n1575), 
        .Y(n503) );
  OAI2BB2XL U1015 ( .B0(n1500), .B1(n1573), .A0N(\gbuff[11][6] ), .A1N(n1575), 
        .Y(n504) );
  OAI2BB2XL U1016 ( .B0(n1498), .B1(n1573), .A0N(\gbuff[11][7] ), .A1N(n1575), 
        .Y(n505) );
  OAI2BB2XL U1017 ( .B0(n1496), .B1(n1573), .A0N(\gbuff[11][8] ), .A1N(n1575), 
        .Y(n506) );
  OAI2BB2XL U1018 ( .B0(n1494), .B1(n1573), .A0N(\gbuff[11][9] ), .A1N(n1575), 
        .Y(n507) );
  OAI2BB2XL U1019 ( .B0(n1492), .B1(n1573), .A0N(\gbuff[11][10] ), .A1N(n1575), 
        .Y(n508) );
  OAI2BB2XL U1020 ( .B0(n1490), .B1(n1573), .A0N(\gbuff[11][11] ), .A1N(n1575), 
        .Y(n509) );
  OAI2BB2XL U1021 ( .B0(n1488), .B1(n1573), .A0N(\gbuff[11][12] ), .A1N(n1575), 
        .Y(n510) );
  OAI2BB2XL U1022 ( .B0(n1486), .B1(n1573), .A0N(\gbuff[11][13] ), .A1N(n1575), 
        .Y(n511) );
  OAI2BB2XL U1023 ( .B0(n1484), .B1(n1574), .A0N(\gbuff[11][14] ), .A1N(n1575), 
        .Y(n512) );
  OAI2BB2XL U1024 ( .B0(n1482), .B1(n1573), .A0N(\gbuff[11][15] ), .A1N(n1574), 
        .Y(n513) );
  OAI2BB2XL U1025 ( .B0(n1480), .B1(n1574), .A0N(\gbuff[11][16] ), .A1N(n1575), 
        .Y(n514) );
  OAI2BB2XL U1026 ( .B0(n1478), .B1(n1573), .A0N(\gbuff[11][17] ), .A1N(n1574), 
        .Y(n515) );
  OAI2BB2XL U1027 ( .B0(n1476), .B1(n1574), .A0N(\gbuff[11][18] ), .A1N(n1574), 
        .Y(n516) );
  OAI2BB2XL U1028 ( .B0(n1474), .B1(n1573), .A0N(\gbuff[11][19] ), .A1N(n1574), 
        .Y(n517) );
  OAI2BB2XL U1029 ( .B0(n1472), .B1(n1574), .A0N(\gbuff[11][20] ), .A1N(n1574), 
        .Y(n518) );
  OAI2BB2XL U1030 ( .B0(n1470), .B1(n1573), .A0N(\gbuff[11][21] ), .A1N(n1574), 
        .Y(n519) );
  OAI2BB2XL U1031 ( .B0(n1468), .B1(n1574), .A0N(\gbuff[11][22] ), .A1N(n1575), 
        .Y(n520) );
  OAI2BB2XL U1032 ( .B0(n1466), .B1(n1574), .A0N(\gbuff[11][23] ), .A1N(n1574), 
        .Y(n521) );
  OAI2BB2XL U1033 ( .B0(n1464), .B1(n1573), .A0N(\gbuff[11][24] ), .A1N(n1575), 
        .Y(n522) );
  OAI2BB2XL U1034 ( .B0(n1462), .B1(n1574), .A0N(\gbuff[11][25] ), .A1N(n1575), 
        .Y(n523) );
  OAI2BB2XL U1035 ( .B0(n1460), .B1(n1574), .A0N(\gbuff[11][26] ), .A1N(n1575), 
        .Y(n524) );
  OAI2BB2XL U1036 ( .B0(n1458), .B1(n1574), .A0N(\gbuff[11][27] ), .A1N(n1575), 
        .Y(n525) );
  OAI2BB2XL U1037 ( .B0(n1456), .B1(n1574), .A0N(\gbuff[11][28] ), .A1N(n1575), 
        .Y(n526) );
  OAI2BB2XL U1038 ( .B0(n1454), .B1(n1574), .A0N(\gbuff[11][29] ), .A1N(n1575), 
        .Y(n527) );
  OAI2BB2XL U1039 ( .B0(n1452), .B1(n1574), .A0N(\gbuff[11][30] ), .A1N(n1575), 
        .Y(n528) );
  OAI2BB2XL U1040 ( .B0(n1450), .B1(n1574), .A0N(\gbuff[11][31] ), .A1N(n1573), 
        .Y(n529) );
  OAI2BB2XL U1041 ( .B0(n1512), .B1(n1570), .A0N(\gbuff[12][0] ), .A1N(n1572), 
        .Y(n530) );
  OAI2BB2XL U1042 ( .B0(n1510), .B1(n1570), .A0N(\gbuff[12][1] ), .A1N(n1570), 
        .Y(n531) );
  OAI2BB2XL U1043 ( .B0(n1508), .B1(n1570), .A0N(\gbuff[12][2] ), .A1N(n1570), 
        .Y(n532) );
  OAI2BB2XL U1044 ( .B0(n1506), .B1(n1570), .A0N(\gbuff[12][3] ), .A1N(n1572), 
        .Y(n533) );
  OAI2BB2XL U1045 ( .B0(n1504), .B1(n1570), .A0N(\gbuff[12][4] ), .A1N(n1570), 
        .Y(n534) );
  OAI2BB2XL U1046 ( .B0(n1502), .B1(n1570), .A0N(\gbuff[12][5] ), .A1N(n1572), 
        .Y(n535) );
  OAI2BB2XL U1047 ( .B0(n1500), .B1(n1570), .A0N(\gbuff[12][6] ), .A1N(n1572), 
        .Y(n536) );
  OAI2BB2XL U1048 ( .B0(n1498), .B1(n1570), .A0N(\gbuff[12][7] ), .A1N(n1572), 
        .Y(n537) );
  OAI2BB2XL U1049 ( .B0(n1496), .B1(n1570), .A0N(\gbuff[12][8] ), .A1N(n1572), 
        .Y(n538) );
  OAI2BB2XL U1050 ( .B0(n1494), .B1(n1570), .A0N(\gbuff[12][9] ), .A1N(n1572), 
        .Y(n539) );
  OAI2BB2XL U1051 ( .B0(n1492), .B1(n1570), .A0N(\gbuff[12][10] ), .A1N(n1572), 
        .Y(n540) );
  OAI2BB2XL U1052 ( .B0(n1490), .B1(n1570), .A0N(\gbuff[12][11] ), .A1N(n1572), 
        .Y(n541) );
  OAI2BB2XL U1053 ( .B0(n1488), .B1(n1570), .A0N(\gbuff[12][12] ), .A1N(n1572), 
        .Y(n542) );
  OAI2BB2XL U1054 ( .B0(n1486), .B1(n1571), .A0N(\gbuff[12][13] ), .A1N(n1572), 
        .Y(n543) );
  OAI2BB2XL U1055 ( .B0(n1484), .B1(n1570), .A0N(\gbuff[12][14] ), .A1N(n1572), 
        .Y(n544) );
  OAI2BB2XL U1056 ( .B0(n1482), .B1(n1571), .A0N(\gbuff[12][15] ), .A1N(n1571), 
        .Y(n545) );
  OAI2BB2XL U1057 ( .B0(n1480), .B1(n1570), .A0N(\gbuff[12][16] ), .A1N(n1572), 
        .Y(n546) );
  OAI2BB2XL U1058 ( .B0(n1478), .B1(n1571), .A0N(\gbuff[12][17] ), .A1N(n1571), 
        .Y(n547) );
  OAI2BB2XL U1059 ( .B0(n1476), .B1(n1570), .A0N(\gbuff[12][18] ), .A1N(n1571), 
        .Y(n548) );
  OAI2BB2XL U1060 ( .B0(n1474), .B1(n1571), .A0N(\gbuff[12][19] ), .A1N(n1571), 
        .Y(n549) );
  OAI2BB2XL U1061 ( .B0(n1472), .B1(n1570), .A0N(\gbuff[12][20] ), .A1N(n1571), 
        .Y(n550) );
  OAI2BB2XL U1062 ( .B0(n1470), .B1(n1571), .A0N(\gbuff[12][21] ), .A1N(n1571), 
        .Y(n551) );
  OAI2BB2XL U1063 ( .B0(n1468), .B1(n1570), .A0N(\gbuff[12][22] ), .A1N(n1572), 
        .Y(n552) );
  OAI2BB2XL U1064 ( .B0(n1466), .B1(n1571), .A0N(\gbuff[12][23] ), .A1N(n1571), 
        .Y(n553) );
  OAI2BB2XL U1065 ( .B0(n1464), .B1(n1571), .A0N(\gbuff[12][24] ), .A1N(n1572), 
        .Y(n554) );
  OAI2BB2XL U1066 ( .B0(n1462), .B1(n1571), .A0N(\gbuff[12][25] ), .A1N(n1572), 
        .Y(n555) );
  OAI2BB2XL U1067 ( .B0(n1460), .B1(n1571), .A0N(\gbuff[12][26] ), .A1N(n1572), 
        .Y(n556) );
  OAI2BB2XL U1068 ( .B0(n1458), .B1(n1571), .A0N(\gbuff[12][27] ), .A1N(n1572), 
        .Y(n557) );
  OAI2BB2XL U1069 ( .B0(n1456), .B1(n1571), .A0N(\gbuff[12][28] ), .A1N(n1572), 
        .Y(n558) );
  OAI2BB2XL U1070 ( .B0(n1454), .B1(n1571), .A0N(\gbuff[12][29] ), .A1N(n1572), 
        .Y(n559) );
  OAI2BB2XL U1071 ( .B0(n1452), .B1(n1571), .A0N(\gbuff[12][30] ), .A1N(n1572), 
        .Y(n560) );
  OAI2BB2XL U1072 ( .B0(n1450), .B1(n1571), .A0N(\gbuff[12][31] ), .A1N(n1572), 
        .Y(n561) );
  OAI2BB2XL U1073 ( .B0(n1512), .B1(n1567), .A0N(\gbuff[13][0] ), .A1N(n1569), 
        .Y(n562) );
  OAI2BB2XL U1074 ( .B0(n1510), .B1(n1567), .A0N(\gbuff[13][1] ), .A1N(n14), 
        .Y(n563) );
  OAI2BB2XL U1075 ( .B0(n1508), .B1(n1567), .A0N(\gbuff[13][2] ), .A1N(n1567), 
        .Y(n564) );
  OAI2BB2XL U1076 ( .B0(n1506), .B1(n1567), .A0N(\gbuff[13][3] ), .A1N(n1569), 
        .Y(n565) );
  OAI2BB2XL U1077 ( .B0(n1504), .B1(n1567), .A0N(\gbuff[13][4] ), .A1N(n1569), 
        .Y(n566) );
  OAI2BB2XL U1078 ( .B0(n1502), .B1(n1567), .A0N(\gbuff[13][5] ), .A1N(n1569), 
        .Y(n567) );
  OAI2BB2XL U1079 ( .B0(n1500), .B1(n1567), .A0N(\gbuff[13][6] ), .A1N(n1569), 
        .Y(n568) );
  OAI2BB2XL U1080 ( .B0(n1498), .B1(n1567), .A0N(\gbuff[13][7] ), .A1N(n1569), 
        .Y(n569) );
  OAI2BB2XL U1081 ( .B0(n1496), .B1(n1567), .A0N(\gbuff[13][8] ), .A1N(n1569), 
        .Y(n570) );
  OAI2BB2XL U1082 ( .B0(n1494), .B1(n1567), .A0N(\gbuff[13][9] ), .A1N(n1569), 
        .Y(n571) );
  OAI2BB2XL U1083 ( .B0(n1492), .B1(n1567), .A0N(\gbuff[13][10] ), .A1N(n1569), 
        .Y(n572) );
  OAI2BB2XL U1084 ( .B0(n1490), .B1(n1567), .A0N(\gbuff[13][11] ), .A1N(n1569), 
        .Y(n573) );
  OAI2BB2XL U1085 ( .B0(n1488), .B1(n1567), .A0N(\gbuff[13][12] ), .A1N(n1569), 
        .Y(n574) );
  OAI2BB2XL U1086 ( .B0(n1486), .B1(n1567), .A0N(\gbuff[13][13] ), .A1N(n1569), 
        .Y(n575) );
  OAI2BB2XL U1087 ( .B0(n1484), .B1(n1568), .A0N(\gbuff[13][14] ), .A1N(n1569), 
        .Y(n576) );
  OAI2BB2XL U1088 ( .B0(n1482), .B1(n1567), .A0N(\gbuff[13][15] ), .A1N(n1568), 
        .Y(n577) );
  OAI2BB2XL U1089 ( .B0(n1480), .B1(n1568), .A0N(\gbuff[13][16] ), .A1N(n1569), 
        .Y(n578) );
  OAI2BB2XL U1090 ( .B0(n1478), .B1(n1567), .A0N(\gbuff[13][17] ), .A1N(n1568), 
        .Y(n579) );
  OAI2BB2XL U1091 ( .B0(n1476), .B1(n1568), .A0N(\gbuff[13][18] ), .A1N(n1568), 
        .Y(n580) );
  OAI2BB2XL U1092 ( .B0(n1474), .B1(n1567), .A0N(\gbuff[13][19] ), .A1N(n1568), 
        .Y(n581) );
  OAI2BB2XL U1093 ( .B0(n1472), .B1(n1568), .A0N(\gbuff[13][20] ), .A1N(n1568), 
        .Y(n582) );
  OAI2BB2XL U1094 ( .B0(n1470), .B1(n1567), .A0N(\gbuff[13][21] ), .A1N(n1568), 
        .Y(n583) );
  OAI2BB2XL U1095 ( .B0(n1468), .B1(n1568), .A0N(\gbuff[13][22] ), .A1N(n1569), 
        .Y(n584) );
  OAI2BB2XL U1096 ( .B0(n1466), .B1(n1568), .A0N(\gbuff[13][23] ), .A1N(n1568), 
        .Y(n585) );
  OAI2BB2XL U1097 ( .B0(n1464), .B1(n14), .A0N(\gbuff[13][24] ), .A1N(n1569), 
        .Y(n586) );
  OAI2BB2XL U1098 ( .B0(n1462), .B1(n1568), .A0N(\gbuff[13][25] ), .A1N(n1569), 
        .Y(n587) );
  OAI2BB2XL U1099 ( .B0(n1460), .B1(n1568), .A0N(\gbuff[13][26] ), .A1N(n1569), 
        .Y(n588) );
  OAI2BB2XL U1100 ( .B0(n1458), .B1(n1568), .A0N(\gbuff[13][27] ), .A1N(n1569), 
        .Y(n589) );
  OAI2BB2XL U1101 ( .B0(n1456), .B1(n1568), .A0N(\gbuff[13][28] ), .A1N(n1569), 
        .Y(n590) );
  OAI2BB2XL U1102 ( .B0(n1454), .B1(n1568), .A0N(\gbuff[13][29] ), .A1N(n1569), 
        .Y(n591) );
  OAI2BB2XL U1103 ( .B0(n1452), .B1(n1568), .A0N(\gbuff[13][30] ), .A1N(n1569), 
        .Y(n592) );
  OAI2BB2XL U1104 ( .B0(n1450), .B1(n1568), .A0N(\gbuff[13][31] ), .A1N(n1567), 
        .Y(n593) );
  OAI2BB2XL U1105 ( .B0(n1512), .B1(n1564), .A0N(\gbuff[14][0] ), .A1N(n1566), 
        .Y(n594) );
  OAI2BB2XL U1106 ( .B0(n1510), .B1(n1564), .A0N(\gbuff[14][1] ), .A1N(n15), 
        .Y(n595) );
  OAI2BB2XL U1107 ( .B0(n1508), .B1(n1564), .A0N(\gbuff[14][2] ), .A1N(n1564), 
        .Y(n596) );
  OAI2BB2XL U1108 ( .B0(n1506), .B1(n1564), .A0N(\gbuff[14][3] ), .A1N(n1566), 
        .Y(n597) );
  OAI2BB2XL U1109 ( .B0(n1504), .B1(n1564), .A0N(\gbuff[14][4] ), .A1N(n1566), 
        .Y(n598) );
  OAI2BB2XL U1110 ( .B0(n1502), .B1(n1564), .A0N(\gbuff[14][5] ), .A1N(n1566), 
        .Y(n599) );
  OAI2BB2XL U1111 ( .B0(n1500), .B1(n1564), .A0N(\gbuff[14][6] ), .A1N(n1566), 
        .Y(n600) );
  OAI2BB2XL U1112 ( .B0(n1498), .B1(n1564), .A0N(\gbuff[14][7] ), .A1N(n1566), 
        .Y(n601) );
  OAI2BB2XL U1113 ( .B0(n1496), .B1(n1564), .A0N(\gbuff[14][8] ), .A1N(n1566), 
        .Y(n602) );
  OAI2BB2XL U1114 ( .B0(n1494), .B1(n1564), .A0N(\gbuff[14][9] ), .A1N(n1566), 
        .Y(n603) );
  OAI2BB2XL U1115 ( .B0(n1492), .B1(n1564), .A0N(\gbuff[14][10] ), .A1N(n1566), 
        .Y(n604) );
  OAI2BB2XL U1116 ( .B0(n1490), .B1(n1564), .A0N(\gbuff[14][11] ), .A1N(n1566), 
        .Y(n605) );
  OAI2BB2XL U1117 ( .B0(n1488), .B1(n1564), .A0N(\gbuff[14][12] ), .A1N(n1566), 
        .Y(n606) );
  OAI2BB2XL U1118 ( .B0(n1486), .B1(n1564), .A0N(\gbuff[14][13] ), .A1N(n1566), 
        .Y(n607) );
  OAI2BB2XL U1119 ( .B0(n1484), .B1(n1565), .A0N(\gbuff[14][14] ), .A1N(n1566), 
        .Y(n608) );
  OAI2BB2XL U1120 ( .B0(n1482), .B1(n1564), .A0N(\gbuff[14][15] ), .A1N(n1565), 
        .Y(n609) );
  OAI2BB2XL U1121 ( .B0(n1480), .B1(n1565), .A0N(\gbuff[14][16] ), .A1N(n1566), 
        .Y(n610) );
  OAI2BB2XL U1122 ( .B0(n1478), .B1(n1564), .A0N(\gbuff[14][17] ), .A1N(n1565), 
        .Y(n611) );
  OAI2BB2XL U1123 ( .B0(n1476), .B1(n1565), .A0N(\gbuff[14][18] ), .A1N(n1565), 
        .Y(n612) );
  OAI2BB2XL U1124 ( .B0(n1474), .B1(n1564), .A0N(\gbuff[14][19] ), .A1N(n1565), 
        .Y(n613) );
  OAI2BB2XL U1125 ( .B0(n1472), .B1(n1565), .A0N(\gbuff[14][20] ), .A1N(n1565), 
        .Y(n614) );
  OAI2BB2XL U1126 ( .B0(n1470), .B1(n1564), .A0N(\gbuff[14][21] ), .A1N(n1565), 
        .Y(n615) );
  OAI2BB2XL U1127 ( .B0(n1468), .B1(n1565), .A0N(\gbuff[14][22] ), .A1N(n1566), 
        .Y(n616) );
  OAI2BB2XL U1128 ( .B0(n1466), .B1(n1565), .A0N(\gbuff[14][23] ), .A1N(n1565), 
        .Y(n617) );
  OAI2BB2XL U1129 ( .B0(n1464), .B1(n15), .A0N(\gbuff[14][24] ), .A1N(n1566), 
        .Y(n618) );
  OAI2BB2XL U1130 ( .B0(n1462), .B1(n1565), .A0N(\gbuff[14][25] ), .A1N(n1566), 
        .Y(n619) );
  OAI2BB2XL U1131 ( .B0(n1460), .B1(n1565), .A0N(\gbuff[14][26] ), .A1N(n1566), 
        .Y(n620) );
  OAI2BB2XL U1132 ( .B0(n1458), .B1(n1565), .A0N(\gbuff[14][27] ), .A1N(n1566), 
        .Y(n621) );
  OAI2BB2XL U1133 ( .B0(n1456), .B1(n1565), .A0N(\gbuff[14][28] ), .A1N(n1566), 
        .Y(n622) );
  OAI2BB2XL U1134 ( .B0(n1454), .B1(n1565), .A0N(\gbuff[14][29] ), .A1N(n1566), 
        .Y(n623) );
  OAI2BB2XL U1135 ( .B0(n1452), .B1(n1565), .A0N(\gbuff[14][30] ), .A1N(n1566), 
        .Y(n624) );
  OAI2BB2XL U1136 ( .B0(n1450), .B1(n1565), .A0N(\gbuff[14][31] ), .A1N(n1564), 
        .Y(n625) );
  OAI2BB2XL U1137 ( .B0(n1512), .B1(n1561), .A0N(\gbuff[15][0] ), .A1N(n1563), 
        .Y(n626) );
  OAI2BB2XL U1138 ( .B0(n1510), .B1(n1561), .A0N(\gbuff[15][1] ), .A1N(n16), 
        .Y(n627) );
  OAI2BB2XL U1139 ( .B0(n1508), .B1(n1561), .A0N(\gbuff[15][2] ), .A1N(n1561), 
        .Y(n628) );
  OAI2BB2XL U1140 ( .B0(n1506), .B1(n1561), .A0N(\gbuff[15][3] ), .A1N(n1563), 
        .Y(n629) );
  OAI2BB2XL U1141 ( .B0(n1504), .B1(n1561), .A0N(\gbuff[15][4] ), .A1N(n1563), 
        .Y(n630) );
  OAI2BB2XL U1142 ( .B0(n1502), .B1(n1561), .A0N(\gbuff[15][5] ), .A1N(n1563), 
        .Y(n631) );
  OAI2BB2XL U1143 ( .B0(n1500), .B1(n1561), .A0N(\gbuff[15][6] ), .A1N(n1563), 
        .Y(n632) );
  OAI2BB2XL U1144 ( .B0(n1498), .B1(n1561), .A0N(\gbuff[15][7] ), .A1N(n1563), 
        .Y(n633) );
  OAI2BB2XL U1145 ( .B0(n1496), .B1(n1561), .A0N(\gbuff[15][8] ), .A1N(n1563), 
        .Y(n634) );
  OAI2BB2XL U1146 ( .B0(n1494), .B1(n1561), .A0N(\gbuff[15][9] ), .A1N(n1563), 
        .Y(n635) );
  OAI2BB2XL U1147 ( .B0(n1492), .B1(n1561), .A0N(\gbuff[15][10] ), .A1N(n1563), 
        .Y(n636) );
  OAI2BB2XL U1148 ( .B0(n1490), .B1(n1561), .A0N(\gbuff[15][11] ), .A1N(n1563), 
        .Y(n637) );
  OAI2BB2XL U1149 ( .B0(n1488), .B1(n1561), .A0N(\gbuff[15][12] ), .A1N(n1563), 
        .Y(n638) );
  OAI2BB2XL U1150 ( .B0(n1486), .B1(n1561), .A0N(\gbuff[15][13] ), .A1N(n1563), 
        .Y(n639) );
  OAI2BB2XL U1151 ( .B0(n1484), .B1(n1562), .A0N(\gbuff[15][14] ), .A1N(n1563), 
        .Y(n640) );
  OAI2BB2XL U1152 ( .B0(n1482), .B1(n1561), .A0N(\gbuff[15][15] ), .A1N(n1562), 
        .Y(n641) );
  OAI2BB2XL U1153 ( .B0(n1480), .B1(n1562), .A0N(\gbuff[15][16] ), .A1N(n1563), 
        .Y(n642) );
  OAI2BB2XL U1154 ( .B0(n1478), .B1(n1561), .A0N(\gbuff[15][17] ), .A1N(n1562), 
        .Y(n643) );
  OAI2BB2XL U1155 ( .B0(n1476), .B1(n1562), .A0N(\gbuff[15][18] ), .A1N(n1562), 
        .Y(n644) );
  OAI2BB2XL U1156 ( .B0(n1474), .B1(n1561), .A0N(\gbuff[15][19] ), .A1N(n1562), 
        .Y(n645) );
  OAI2BB2XL U1157 ( .B0(n1472), .B1(n1562), .A0N(\gbuff[15][20] ), .A1N(n1562), 
        .Y(n646) );
  OAI2BB2XL U1158 ( .B0(n1470), .B1(n1561), .A0N(\gbuff[15][21] ), .A1N(n1562), 
        .Y(n647) );
  OAI2BB2XL U1159 ( .B0(n1468), .B1(n1562), .A0N(\gbuff[15][22] ), .A1N(n1563), 
        .Y(n648) );
  OAI2BB2XL U1160 ( .B0(n1466), .B1(n1562), .A0N(\gbuff[15][23] ), .A1N(n1562), 
        .Y(n649) );
  OAI2BB2XL U1161 ( .B0(n1464), .B1(n16), .A0N(\gbuff[15][24] ), .A1N(n1563), 
        .Y(n650) );
  OAI2BB2XL U1162 ( .B0(n1462), .B1(n1562), .A0N(\gbuff[15][25] ), .A1N(n1563), 
        .Y(n651) );
  OAI2BB2XL U1163 ( .B0(n1460), .B1(n1562), .A0N(\gbuff[15][26] ), .A1N(n1563), 
        .Y(n652) );
  OAI2BB2XL U1164 ( .B0(n1458), .B1(n1562), .A0N(\gbuff[15][27] ), .A1N(n1563), 
        .Y(n653) );
  OAI2BB2XL U1165 ( .B0(n1456), .B1(n1562), .A0N(\gbuff[15][28] ), .A1N(n1563), 
        .Y(n654) );
  OAI2BB2XL U1166 ( .B0(n1454), .B1(n1562), .A0N(\gbuff[15][29] ), .A1N(n1563), 
        .Y(n655) );
  OAI2BB2XL U1167 ( .B0(n1452), .B1(n1562), .A0N(\gbuff[15][30] ), .A1N(n1563), 
        .Y(n656) );
  OAI2BB2XL U1168 ( .B0(n1450), .B1(n1562), .A0N(\gbuff[15][31] ), .A1N(n1561), 
        .Y(n657) );
  OAI2BB2XL U1169 ( .B0(n1512), .B1(n1558), .A0N(\gbuff[16][0] ), .A1N(n1560), 
        .Y(n658) );
  OAI2BB2XL U1170 ( .B0(n1510), .B1(n1558), .A0N(\gbuff[16][1] ), .A1N(n1559), 
        .Y(n659) );
  OAI2BB2XL U1171 ( .B0(n1508), .B1(n1558), .A0N(\gbuff[16][2] ), .A1N(n1558), 
        .Y(n660) );
  OAI2BB2XL U1172 ( .B0(n1506), .B1(n1558), .A0N(\gbuff[16][3] ), .A1N(n1560), 
        .Y(n661) );
  OAI2BB2XL U1173 ( .B0(n1504), .B1(n1558), .A0N(\gbuff[16][4] ), .A1N(n1560), 
        .Y(n662) );
  OAI2BB2XL U1174 ( .B0(n1502), .B1(n1558), .A0N(\gbuff[16][5] ), .A1N(n1560), 
        .Y(n663) );
  OAI2BB2XL U1175 ( .B0(n1500), .B1(n1558), .A0N(\gbuff[16][6] ), .A1N(n1560), 
        .Y(n664) );
  OAI2BB2XL U1176 ( .B0(n1498), .B1(n1558), .A0N(\gbuff[16][7] ), .A1N(n1560), 
        .Y(n665) );
  OAI2BB2XL U1177 ( .B0(n1496), .B1(n1558), .A0N(\gbuff[16][8] ), .A1N(n1560), 
        .Y(n666) );
  OAI2BB2XL U1178 ( .B0(n1494), .B1(n1558), .A0N(\gbuff[16][9] ), .A1N(n1560), 
        .Y(n667) );
  OAI2BB2XL U1179 ( .B0(n1492), .B1(n1558), .A0N(\gbuff[16][10] ), .A1N(n1560), 
        .Y(n668) );
  OAI2BB2XL U1180 ( .B0(n1490), .B1(n1558), .A0N(\gbuff[16][11] ), .A1N(n1560), 
        .Y(n669) );
  OAI2BB2XL U1181 ( .B0(n1488), .B1(n1558), .A0N(\gbuff[16][12] ), .A1N(n1560), 
        .Y(n670) );
  OAI2BB2XL U1182 ( .B0(n1486), .B1(n1558), .A0N(\gbuff[16][13] ), .A1N(n1560), 
        .Y(n671) );
  OAI2BB2XL U1183 ( .B0(n1484), .B1(n1559), .A0N(\gbuff[16][14] ), .A1N(n1560), 
        .Y(n672) );
  OAI2BB2XL U1184 ( .B0(n1482), .B1(n1558), .A0N(\gbuff[16][15] ), .A1N(n1559), 
        .Y(n673) );
  OAI2BB2XL U1185 ( .B0(n1480), .B1(n1559), .A0N(\gbuff[16][16] ), .A1N(n1560), 
        .Y(n674) );
  OAI2BB2XL U1186 ( .B0(n1478), .B1(n1558), .A0N(\gbuff[16][17] ), .A1N(n1559), 
        .Y(n675) );
  OAI2BB2XL U1187 ( .B0(n1476), .B1(n1559), .A0N(\gbuff[16][18] ), .A1N(n1559), 
        .Y(n676) );
  OAI2BB2XL U1188 ( .B0(n1474), .B1(n1558), .A0N(\gbuff[16][19] ), .A1N(n1559), 
        .Y(n677) );
  OAI2BB2XL U1189 ( .B0(n1472), .B1(n1559), .A0N(\gbuff[16][20] ), .A1N(n1559), 
        .Y(n678) );
  OAI2BB2XL U1190 ( .B0(n1470), .B1(n1558), .A0N(\gbuff[16][21] ), .A1N(n1559), 
        .Y(n679) );
  OAI2BB2XL U1191 ( .B0(n1468), .B1(n1559), .A0N(\gbuff[16][22] ), .A1N(n1560), 
        .Y(n680) );
  OAI2BB2XL U1192 ( .B0(n1466), .B1(n1559), .A0N(\gbuff[16][23] ), .A1N(n1559), 
        .Y(n681) );
  OAI2BB2XL U1193 ( .B0(n1464), .B1(n1558), .A0N(\gbuff[16][24] ), .A1N(n1560), 
        .Y(n682) );
  OAI2BB2XL U1194 ( .B0(n1462), .B1(n1559), .A0N(\gbuff[16][25] ), .A1N(n1560), 
        .Y(n683) );
  OAI2BB2XL U1195 ( .B0(n1460), .B1(n1559), .A0N(\gbuff[16][26] ), .A1N(n1560), 
        .Y(n684) );
  OAI2BB2XL U1196 ( .B0(n1458), .B1(n1559), .A0N(\gbuff[16][27] ), .A1N(n1560), 
        .Y(n685) );
  OAI2BB2XL U1197 ( .B0(n1456), .B1(n1559), .A0N(\gbuff[16][28] ), .A1N(n1560), 
        .Y(n686) );
  OAI2BB2XL U1198 ( .B0(n1454), .B1(n1559), .A0N(\gbuff[16][29] ), .A1N(n1560), 
        .Y(n687) );
  OAI2BB2XL U1199 ( .B0(n1452), .B1(n1559), .A0N(\gbuff[16][30] ), .A1N(n1560), 
        .Y(n688) );
  OAI2BB2XL U1200 ( .B0(n1450), .B1(n1559), .A0N(\gbuff[16][31] ), .A1N(n1558), 
        .Y(n689) );
  OAI2BB2XL U1201 ( .B0(n1512), .B1(n1555), .A0N(\gbuff[17][0] ), .A1N(n1557), 
        .Y(n690) );
  OAI2BB2XL U1202 ( .B0(n1510), .B1(n1555), .A0N(\gbuff[17][1] ), .A1N(n1556), 
        .Y(n691) );
  OAI2BB2XL U1203 ( .B0(n1508), .B1(n1555), .A0N(\gbuff[17][2] ), .A1N(n1555), 
        .Y(n692) );
  OAI2BB2XL U1204 ( .B0(n1506), .B1(n1555), .A0N(\gbuff[17][3] ), .A1N(n1557), 
        .Y(n693) );
  OAI2BB2XL U1205 ( .B0(n1504), .B1(n1555), .A0N(\gbuff[17][4] ), .A1N(n1557), 
        .Y(n694) );
  OAI2BB2XL U1206 ( .B0(n1502), .B1(n1555), .A0N(\gbuff[17][5] ), .A1N(n1557), 
        .Y(n695) );
  OAI2BB2XL U1207 ( .B0(n1500), .B1(n1555), .A0N(\gbuff[17][6] ), .A1N(n1557), 
        .Y(n696) );
  OAI2BB2XL U1208 ( .B0(n1498), .B1(n1555), .A0N(\gbuff[17][7] ), .A1N(n1557), 
        .Y(n697) );
  OAI2BB2XL U1209 ( .B0(n1496), .B1(n1555), .A0N(\gbuff[17][8] ), .A1N(n1557), 
        .Y(n698) );
  OAI2BB2XL U1210 ( .B0(n1494), .B1(n1555), .A0N(\gbuff[17][9] ), .A1N(n1557), 
        .Y(n699) );
  OAI2BB2XL U1211 ( .B0(n1492), .B1(n1555), .A0N(\gbuff[17][10] ), .A1N(n1557), 
        .Y(n700) );
  OAI2BB2XL U1212 ( .B0(n1490), .B1(n1555), .A0N(\gbuff[17][11] ), .A1N(n1557), 
        .Y(n701) );
  OAI2BB2XL U1213 ( .B0(n1488), .B1(n1555), .A0N(\gbuff[17][12] ), .A1N(n1557), 
        .Y(n702) );
  OAI2BB2XL U1214 ( .B0(n1486), .B1(n1555), .A0N(\gbuff[17][13] ), .A1N(n1557), 
        .Y(n703) );
  OAI2BB2XL U1215 ( .B0(n1484), .B1(n1556), .A0N(\gbuff[17][14] ), .A1N(n1557), 
        .Y(n704) );
  OAI2BB2XL U1216 ( .B0(n1482), .B1(n1555), .A0N(\gbuff[17][15] ), .A1N(n1556), 
        .Y(n705) );
  OAI2BB2XL U1217 ( .B0(n1480), .B1(n1556), .A0N(\gbuff[17][16] ), .A1N(n1557), 
        .Y(n706) );
  OAI2BB2XL U1218 ( .B0(n1478), .B1(n1555), .A0N(\gbuff[17][17] ), .A1N(n1556), 
        .Y(n707) );
  OAI2BB2XL U1219 ( .B0(n1476), .B1(n1556), .A0N(\gbuff[17][18] ), .A1N(n1556), 
        .Y(n708) );
  OAI2BB2XL U1220 ( .B0(n1474), .B1(n1555), .A0N(\gbuff[17][19] ), .A1N(n1556), 
        .Y(n709) );
  OAI2BB2XL U1221 ( .B0(n1472), .B1(n1556), .A0N(\gbuff[17][20] ), .A1N(n1556), 
        .Y(n710) );
  OAI2BB2XL U1222 ( .B0(n1470), .B1(n1555), .A0N(\gbuff[17][21] ), .A1N(n1556), 
        .Y(n711) );
  OAI2BB2XL U1223 ( .B0(n1468), .B1(n1556), .A0N(\gbuff[17][22] ), .A1N(n1557), 
        .Y(n712) );
  OAI2BB2XL U1224 ( .B0(n1466), .B1(n1556), .A0N(\gbuff[17][23] ), .A1N(n1556), 
        .Y(n713) );
  OAI2BB2XL U1225 ( .B0(n1464), .B1(n1555), .A0N(\gbuff[17][24] ), .A1N(n1557), 
        .Y(n714) );
  OAI2BB2XL U1226 ( .B0(n1462), .B1(n1556), .A0N(\gbuff[17][25] ), .A1N(n1557), 
        .Y(n715) );
  OAI2BB2XL U1227 ( .B0(n1460), .B1(n1556), .A0N(\gbuff[17][26] ), .A1N(n1557), 
        .Y(n716) );
  OAI2BB2XL U1228 ( .B0(n1458), .B1(n1556), .A0N(\gbuff[17][27] ), .A1N(n1557), 
        .Y(n717) );
  OAI2BB2XL U1229 ( .B0(n1456), .B1(n1556), .A0N(\gbuff[17][28] ), .A1N(n1557), 
        .Y(n718) );
  OAI2BB2XL U1230 ( .B0(n1454), .B1(n1556), .A0N(\gbuff[17][29] ), .A1N(n1557), 
        .Y(n719) );
  OAI2BB2XL U1231 ( .B0(n1452), .B1(n1556), .A0N(\gbuff[17][30] ), .A1N(n1557), 
        .Y(n720) );
  OAI2BB2XL U1232 ( .B0(n1450), .B1(n1556), .A0N(\gbuff[17][31] ), .A1N(n1555), 
        .Y(n721) );
  OAI2BB2XL U1233 ( .B0(n1512), .B1(n1552), .A0N(\gbuff[18][0] ), .A1N(n1554), 
        .Y(n722) );
  OAI2BB2XL U1234 ( .B0(n1510), .B1(n1552), .A0N(\gbuff[18][1] ), .A1N(n1553), 
        .Y(n723) );
  OAI2BB2XL U1235 ( .B0(n1508), .B1(n1552), .A0N(\gbuff[18][2] ), .A1N(n1552), 
        .Y(n724) );
  OAI2BB2XL U1236 ( .B0(n1506), .B1(n1552), .A0N(\gbuff[18][3] ), .A1N(n1554), 
        .Y(n725) );
  OAI2BB2XL U1237 ( .B0(n1504), .B1(n1552), .A0N(\gbuff[18][4] ), .A1N(n1554), 
        .Y(n726) );
  OAI2BB2XL U1238 ( .B0(n1502), .B1(n1552), .A0N(\gbuff[18][5] ), .A1N(n1554), 
        .Y(n727) );
  OAI2BB2XL U1239 ( .B0(n1500), .B1(n1552), .A0N(\gbuff[18][6] ), .A1N(n1554), 
        .Y(n728) );
  OAI2BB2XL U1240 ( .B0(n1498), .B1(n1552), .A0N(\gbuff[18][7] ), .A1N(n1554), 
        .Y(n729) );
  OAI2BB2XL U1241 ( .B0(n1496), .B1(n1552), .A0N(\gbuff[18][8] ), .A1N(n1554), 
        .Y(n730) );
  OAI2BB2XL U1242 ( .B0(n1494), .B1(n1552), .A0N(\gbuff[18][9] ), .A1N(n1554), 
        .Y(n731) );
  OAI2BB2XL U1243 ( .B0(n1492), .B1(n1552), .A0N(\gbuff[18][10] ), .A1N(n1554), 
        .Y(n732) );
  OAI2BB2XL U1244 ( .B0(n1490), .B1(n1552), .A0N(\gbuff[18][11] ), .A1N(n1554), 
        .Y(n733) );
  OAI2BB2XL U1245 ( .B0(n1488), .B1(n1552), .A0N(\gbuff[18][12] ), .A1N(n1554), 
        .Y(n734) );
  OAI2BB2XL U1246 ( .B0(n1486), .B1(n1552), .A0N(\gbuff[18][13] ), .A1N(n1554), 
        .Y(n735) );
  OAI2BB2XL U1247 ( .B0(n1484), .B1(n1553), .A0N(\gbuff[18][14] ), .A1N(n1554), 
        .Y(n736) );
  OAI2BB2XL U1248 ( .B0(n1482), .B1(n1552), .A0N(\gbuff[18][15] ), .A1N(n1553), 
        .Y(n737) );
  OAI2BB2XL U1249 ( .B0(n1480), .B1(n1553), .A0N(\gbuff[18][16] ), .A1N(n1554), 
        .Y(n738) );
  OAI2BB2XL U1250 ( .B0(n1478), .B1(n1552), .A0N(\gbuff[18][17] ), .A1N(n1553), 
        .Y(n739) );
  OAI2BB2XL U1251 ( .B0(n1476), .B1(n1553), .A0N(\gbuff[18][18] ), .A1N(n1553), 
        .Y(n740) );
  OAI2BB2XL U1252 ( .B0(n1474), .B1(n1552), .A0N(\gbuff[18][19] ), .A1N(n1553), 
        .Y(n741) );
  OAI2BB2XL U1253 ( .B0(n1472), .B1(n1553), .A0N(\gbuff[18][20] ), .A1N(n1553), 
        .Y(n742) );
  OAI2BB2XL U1254 ( .B0(n1470), .B1(n1552), .A0N(\gbuff[18][21] ), .A1N(n1553), 
        .Y(n743) );
  OAI2BB2XL U1255 ( .B0(n1468), .B1(n1553), .A0N(\gbuff[18][22] ), .A1N(n1554), 
        .Y(n744) );
  OAI2BB2XL U1256 ( .B0(n1466), .B1(n1553), .A0N(\gbuff[18][23] ), .A1N(n1553), 
        .Y(n745) );
  OAI2BB2XL U1257 ( .B0(n1464), .B1(n1552), .A0N(\gbuff[18][24] ), .A1N(n1554), 
        .Y(n746) );
  OAI2BB2XL U1258 ( .B0(n1462), .B1(n1553), .A0N(\gbuff[18][25] ), .A1N(n1554), 
        .Y(n747) );
  OAI2BB2XL U1259 ( .B0(n1460), .B1(n1553), .A0N(\gbuff[18][26] ), .A1N(n1554), 
        .Y(n748) );
  OAI2BB2XL U1260 ( .B0(n1458), .B1(n1553), .A0N(\gbuff[18][27] ), .A1N(n1554), 
        .Y(n749) );
  OAI2BB2XL U1261 ( .B0(n1456), .B1(n1553), .A0N(\gbuff[18][28] ), .A1N(n1554), 
        .Y(n750) );
  OAI2BB2XL U1262 ( .B0(n1454), .B1(n1553), .A0N(\gbuff[18][29] ), .A1N(n1554), 
        .Y(n751) );
  OAI2BB2XL U1263 ( .B0(n1452), .B1(n1553), .A0N(\gbuff[18][30] ), .A1N(n1554), 
        .Y(n752) );
  OAI2BB2XL U1264 ( .B0(n1450), .B1(n1553), .A0N(\gbuff[18][31] ), .A1N(n1552), 
        .Y(n753) );
  OAI2BB2XL U1265 ( .B0(n1512), .B1(n1549), .A0N(\gbuff[19][0] ), .A1N(n1551), 
        .Y(n754) );
  OAI2BB2XL U1266 ( .B0(n1510), .B1(n1549), .A0N(\gbuff[19][1] ), .A1N(n1550), 
        .Y(n755) );
  OAI2BB2XL U1267 ( .B0(n1508), .B1(n1549), .A0N(\gbuff[19][2] ), .A1N(n1549), 
        .Y(n756) );
  OAI2BB2XL U1268 ( .B0(n1506), .B1(n1549), .A0N(\gbuff[19][3] ), .A1N(n1551), 
        .Y(n757) );
  OAI2BB2XL U1269 ( .B0(n1504), .B1(n1549), .A0N(\gbuff[19][4] ), .A1N(n1551), 
        .Y(n758) );
  OAI2BB2XL U1270 ( .B0(n1502), .B1(n1549), .A0N(\gbuff[19][5] ), .A1N(n1551), 
        .Y(n759) );
  OAI2BB2XL U1271 ( .B0(n1500), .B1(n1549), .A0N(\gbuff[19][6] ), .A1N(n1551), 
        .Y(n760) );
  OAI2BB2XL U1272 ( .B0(n1498), .B1(n1549), .A0N(\gbuff[19][7] ), .A1N(n1551), 
        .Y(n761) );
  OAI2BB2XL U1273 ( .B0(n1496), .B1(n1549), .A0N(\gbuff[19][8] ), .A1N(n1551), 
        .Y(n762) );
  OAI2BB2XL U1274 ( .B0(n1494), .B1(n1549), .A0N(\gbuff[19][9] ), .A1N(n1551), 
        .Y(n763) );
  OAI2BB2XL U1275 ( .B0(n1492), .B1(n1549), .A0N(\gbuff[19][10] ), .A1N(n1551), 
        .Y(n764) );
  OAI2BB2XL U1276 ( .B0(n1490), .B1(n1549), .A0N(\gbuff[19][11] ), .A1N(n1551), 
        .Y(n765) );
  OAI2BB2XL U1277 ( .B0(n1488), .B1(n1549), .A0N(\gbuff[19][12] ), .A1N(n1551), 
        .Y(n766) );
  OAI2BB2XL U1278 ( .B0(n1486), .B1(n1549), .A0N(\gbuff[19][13] ), .A1N(n1551), 
        .Y(n767) );
  OAI2BB2XL U1279 ( .B0(n1484), .B1(n1550), .A0N(\gbuff[19][14] ), .A1N(n1551), 
        .Y(n768) );
  OAI2BB2XL U1280 ( .B0(n1482), .B1(n1549), .A0N(\gbuff[19][15] ), .A1N(n1550), 
        .Y(n769) );
  OAI2BB2XL U1281 ( .B0(n1480), .B1(n1550), .A0N(\gbuff[19][16] ), .A1N(n1551), 
        .Y(n770) );
  OAI2BB2XL U1282 ( .B0(n1478), .B1(n1549), .A0N(\gbuff[19][17] ), .A1N(n1550), 
        .Y(n771) );
  OAI2BB2XL U1283 ( .B0(n1476), .B1(n1550), .A0N(\gbuff[19][18] ), .A1N(n1550), 
        .Y(n772) );
  OAI2BB2XL U1284 ( .B0(n1474), .B1(n1549), .A0N(\gbuff[19][19] ), .A1N(n1550), 
        .Y(n773) );
  OAI2BB2XL U1285 ( .B0(n1472), .B1(n1550), .A0N(\gbuff[19][20] ), .A1N(n1550), 
        .Y(n774) );
  OAI2BB2XL U1286 ( .B0(n1470), .B1(n1549), .A0N(\gbuff[19][21] ), .A1N(n1550), 
        .Y(n775) );
  OAI2BB2XL U1287 ( .B0(n1468), .B1(n1550), .A0N(\gbuff[19][22] ), .A1N(n1551), 
        .Y(n776) );
  OAI2BB2XL U1288 ( .B0(n1466), .B1(n1550), .A0N(\gbuff[19][23] ), .A1N(n1550), 
        .Y(n777) );
  OAI2BB2XL U1289 ( .B0(n1464), .B1(n1549), .A0N(\gbuff[19][24] ), .A1N(n1551), 
        .Y(n778) );
  OAI2BB2XL U1290 ( .B0(n1462), .B1(n1550), .A0N(\gbuff[19][25] ), .A1N(n1551), 
        .Y(n779) );
  OAI2BB2XL U1291 ( .B0(n1460), .B1(n1550), .A0N(\gbuff[19][26] ), .A1N(n1551), 
        .Y(n780) );
  OAI2BB2XL U1292 ( .B0(n1458), .B1(n1550), .A0N(\gbuff[19][27] ), .A1N(n1551), 
        .Y(n781) );
  OAI2BB2XL U1293 ( .B0(n1456), .B1(n1550), .A0N(\gbuff[19][28] ), .A1N(n1551), 
        .Y(n782) );
  OAI2BB2XL U1294 ( .B0(n1454), .B1(n1550), .A0N(\gbuff[19][29] ), .A1N(n1551), 
        .Y(n783) );
  OAI2BB2XL U1295 ( .B0(n1452), .B1(n1550), .A0N(\gbuff[19][30] ), .A1N(n1551), 
        .Y(n784) );
  OAI2BB2XL U1296 ( .B0(n1450), .B1(n1550), .A0N(\gbuff[19][31] ), .A1N(n1549), 
        .Y(n785) );
  OAI2BB2XL U1297 ( .B0(n1511), .B1(n1547), .A0N(\gbuff[20][0] ), .A1N(n1547), 
        .Y(n786) );
  OAI2BB2XL U1298 ( .B0(n1509), .B1(n1546), .A0N(\gbuff[20][1] ), .A1N(n1546), 
        .Y(n787) );
  OAI2BB2XL U1299 ( .B0(n1507), .B1(n1546), .A0N(\gbuff[20][2] ), .A1N(n1547), 
        .Y(n788) );
  OAI2BB2XL U1300 ( .B0(n1505), .B1(n1546), .A0N(\gbuff[20][3] ), .A1N(n1548), 
        .Y(n789) );
  OAI2BB2XL U1301 ( .B0(n1503), .B1(n1546), .A0N(\gbuff[20][4] ), .A1N(n1546), 
        .Y(n790) );
  OAI2BB2XL U1302 ( .B0(n1501), .B1(n1546), .A0N(\gbuff[20][5] ), .A1N(n1548), 
        .Y(n791) );
  OAI2BB2XL U1303 ( .B0(n1499), .B1(n1546), .A0N(\gbuff[20][6] ), .A1N(n1548), 
        .Y(n792) );
  OAI2BB2XL U1304 ( .B0(n1497), .B1(n1546), .A0N(\gbuff[20][7] ), .A1N(n1548), 
        .Y(n793) );
  OAI2BB2XL U1305 ( .B0(n1495), .B1(n1546), .A0N(\gbuff[20][8] ), .A1N(n1548), 
        .Y(n794) );
  OAI2BB2XL U1306 ( .B0(n1493), .B1(n1546), .A0N(\gbuff[20][9] ), .A1N(n1548), 
        .Y(n795) );
  OAI2BB2XL U1307 ( .B0(n1491), .B1(n1546), .A0N(\gbuff[20][10] ), .A1N(n1548), 
        .Y(n796) );
  OAI2BB2XL U1308 ( .B0(n1489), .B1(n1546), .A0N(\gbuff[20][11] ), .A1N(n1548), 
        .Y(n797) );
  OAI2BB2XL U1309 ( .B0(n1487), .B1(n1546), .A0N(\gbuff[20][12] ), .A1N(n1548), 
        .Y(n798) );
  OAI2BB2XL U1310 ( .B0(n1485), .B1(n1547), .A0N(\gbuff[20][13] ), .A1N(n1548), 
        .Y(n799) );
  OAI2BB2XL U1311 ( .B0(n1483), .B1(n1547), .A0N(\gbuff[20][14] ), .A1N(n1548), 
        .Y(n800) );
  OAI2BB2XL U1312 ( .B0(n1481), .B1(n1547), .A0N(\gbuff[20][15] ), .A1N(n1548), 
        .Y(n801) );
  OAI2BB2XL U1313 ( .B0(n1479), .B1(n1547), .A0N(\gbuff[20][16] ), .A1N(n1548), 
        .Y(n802) );
  OAI2BB2XL U1314 ( .B0(n1477), .B1(n1547), .A0N(\gbuff[20][17] ), .A1N(n1548), 
        .Y(n803) );
  OAI2BB2XL U1315 ( .B0(n1475), .B1(n1547), .A0N(\gbuff[20][18] ), .A1N(n133), 
        .Y(n804) );
  OAI2BB2XL U1316 ( .B0(n1473), .B1(n1547), .A0N(\gbuff[20][19] ), .A1N(n1546), 
        .Y(n805) );
  OAI2BB2XL U1317 ( .B0(n1471), .B1(n1547), .A0N(\gbuff[20][20] ), .A1N(n1547), 
        .Y(n806) );
  OAI2BB2XL U1318 ( .B0(n1469), .B1(n1547), .A0N(\gbuff[20][21] ), .A1N(n133), 
        .Y(n807) );
  OAI2BB2XL U1319 ( .B0(n1467), .B1(n1547), .A0N(\gbuff[20][22] ), .A1N(n1548), 
        .Y(n808) );
  OAI2BB2XL U1320 ( .B0(n1465), .B1(n1546), .A0N(\gbuff[20][23] ), .A1N(n1548), 
        .Y(n809) );
  OAI2BB2XL U1321 ( .B0(n1463), .B1(n1547), .A0N(\gbuff[20][24] ), .A1N(n1548), 
        .Y(n810) );
  OAI2BB2XL U1322 ( .B0(n1461), .B1(n1547), .A0N(\gbuff[20][25] ), .A1N(n1548), 
        .Y(n811) );
  OAI2BB2XL U1323 ( .B0(n1459), .B1(n1546), .A0N(\gbuff[20][26] ), .A1N(n1548), 
        .Y(n812) );
  OAI2BB2XL U1324 ( .B0(n1457), .B1(n1547), .A0N(\gbuff[20][27] ), .A1N(n1548), 
        .Y(n813) );
  OAI2BB2XL U1325 ( .B0(n1455), .B1(n1546), .A0N(\gbuff[20][28] ), .A1N(n1548), 
        .Y(n814) );
  OAI2BB2XL U1326 ( .B0(n1453), .B1(n1547), .A0N(\gbuff[20][29] ), .A1N(n1548), 
        .Y(n815) );
  OAI2BB2XL U1327 ( .B0(n1451), .B1(n1546), .A0N(\gbuff[20][30] ), .A1N(n1547), 
        .Y(n816) );
  OAI2BB2XL U1328 ( .B0(n1449), .B1(n1547), .A0N(\gbuff[20][31] ), .A1N(n1546), 
        .Y(n817) );
  OAI2BB2XL U1329 ( .B0(n1511), .B1(n1543), .A0N(\gbuff[21][0] ), .A1N(n1545), 
        .Y(n818) );
  OAI2BB2XL U1330 ( .B0(n1509), .B1(n1543), .A0N(\gbuff[21][1] ), .A1N(n134), 
        .Y(n819) );
  OAI2BB2XL U1331 ( .B0(n1507), .B1(n1543), .A0N(\gbuff[21][2] ), .A1N(n1543), 
        .Y(n820) );
  OAI2BB2XL U1332 ( .B0(n1505), .B1(n1543), .A0N(\gbuff[21][3] ), .A1N(n1545), 
        .Y(n821) );
  OAI2BB2XL U1333 ( .B0(n1503), .B1(n1543), .A0N(\gbuff[21][4] ), .A1N(n1545), 
        .Y(n822) );
  OAI2BB2XL U1334 ( .B0(n1501), .B1(n1543), .A0N(\gbuff[21][5] ), .A1N(n1545), 
        .Y(n823) );
  OAI2BB2XL U1335 ( .B0(n1499), .B1(n1543), .A0N(\gbuff[21][6] ), .A1N(n1545), 
        .Y(n824) );
  OAI2BB2XL U1336 ( .B0(n1497), .B1(n1543), .A0N(\gbuff[21][7] ), .A1N(n1545), 
        .Y(n825) );
  OAI2BB2XL U1337 ( .B0(n1495), .B1(n1543), .A0N(\gbuff[21][8] ), .A1N(n1545), 
        .Y(n826) );
  OAI2BB2XL U1338 ( .B0(n1493), .B1(n1543), .A0N(\gbuff[21][9] ), .A1N(n1545), 
        .Y(n827) );
  OAI2BB2XL U1339 ( .B0(n1491), .B1(n1543), .A0N(\gbuff[21][10] ), .A1N(n1545), 
        .Y(n828) );
  OAI2BB2XL U1340 ( .B0(n1489), .B1(n1543), .A0N(\gbuff[21][11] ), .A1N(n1545), 
        .Y(n829) );
  OAI2BB2XL U1341 ( .B0(n1487), .B1(n1543), .A0N(\gbuff[21][12] ), .A1N(n1545), 
        .Y(n830) );
  OAI2BB2XL U1342 ( .B0(n1485), .B1(n1543), .A0N(\gbuff[21][13] ), .A1N(n1545), 
        .Y(n831) );
  OAI2BB2XL U1343 ( .B0(n1483), .B1(n1544), .A0N(\gbuff[21][14] ), .A1N(n1545), 
        .Y(n832) );
  OAI2BB2XL U1344 ( .B0(n1481), .B1(n1543), .A0N(\gbuff[21][15] ), .A1N(n1544), 
        .Y(n833) );
  OAI2BB2XL U1345 ( .B0(n1479), .B1(n1544), .A0N(\gbuff[21][16] ), .A1N(n1545), 
        .Y(n834) );
  OAI2BB2XL U1346 ( .B0(n1477), .B1(n1543), .A0N(\gbuff[21][17] ), .A1N(n1544), 
        .Y(n835) );
  OAI2BB2XL U1347 ( .B0(n1475), .B1(n1544), .A0N(\gbuff[21][18] ), .A1N(n1544), 
        .Y(n836) );
  OAI2BB2XL U1348 ( .B0(n1473), .B1(n1543), .A0N(\gbuff[21][19] ), .A1N(n1544), 
        .Y(n837) );
  OAI2BB2XL U1349 ( .B0(n1471), .B1(n1544), .A0N(\gbuff[21][20] ), .A1N(n1544), 
        .Y(n838) );
  OAI2BB2XL U1350 ( .B0(n1469), .B1(n1543), .A0N(\gbuff[21][21] ), .A1N(n1544), 
        .Y(n839) );
  OAI2BB2XL U1351 ( .B0(n1467), .B1(n1544), .A0N(\gbuff[21][22] ), .A1N(n1545), 
        .Y(n840) );
  OAI2BB2XL U1352 ( .B0(n1465), .B1(n1544), .A0N(\gbuff[21][23] ), .A1N(n1544), 
        .Y(n841) );
  OAI2BB2XL U1353 ( .B0(n1463), .B1(n134), .A0N(\gbuff[21][24] ), .A1N(n1545), 
        .Y(n842) );
  OAI2BB2XL U1354 ( .B0(n1461), .B1(n1544), .A0N(\gbuff[21][25] ), .A1N(n1545), 
        .Y(n843) );
  OAI2BB2XL U1355 ( .B0(n1459), .B1(n1544), .A0N(\gbuff[21][26] ), .A1N(n1545), 
        .Y(n844) );
  OAI2BB2XL U1356 ( .B0(n1457), .B1(n1544), .A0N(\gbuff[21][27] ), .A1N(n1545), 
        .Y(n845) );
  OAI2BB2XL U1357 ( .B0(n1455), .B1(n1544), .A0N(\gbuff[21][28] ), .A1N(n1545), 
        .Y(n846) );
  OAI2BB2XL U1358 ( .B0(n1453), .B1(n1544), .A0N(\gbuff[21][29] ), .A1N(n1545), 
        .Y(n847) );
  OAI2BB2XL U1359 ( .B0(n1451), .B1(n1544), .A0N(\gbuff[21][30] ), .A1N(n1545), 
        .Y(n848) );
  OAI2BB2XL U1360 ( .B0(n1449), .B1(n1544), .A0N(\gbuff[21][31] ), .A1N(n1543), 
        .Y(n849) );
  OAI2BB2XL U1361 ( .B0(n1511), .B1(n1540), .A0N(\gbuff[22][0] ), .A1N(n1542), 
        .Y(n850) );
  OAI2BB2XL U1362 ( .B0(n1509), .B1(n1540), .A0N(\gbuff[22][1] ), .A1N(n135), 
        .Y(n851) );
  OAI2BB2XL U1363 ( .B0(n1507), .B1(n1540), .A0N(\gbuff[22][2] ), .A1N(n1540), 
        .Y(n852) );
  OAI2BB2XL U1364 ( .B0(n1505), .B1(n1540), .A0N(\gbuff[22][3] ), .A1N(n1542), 
        .Y(n853) );
  OAI2BB2XL U1365 ( .B0(n1503), .B1(n1540), .A0N(\gbuff[22][4] ), .A1N(n1542), 
        .Y(n854) );
  OAI2BB2XL U1366 ( .B0(n1501), .B1(n1540), .A0N(\gbuff[22][5] ), .A1N(n1542), 
        .Y(n855) );
  OAI2BB2XL U1367 ( .B0(n1499), .B1(n1540), .A0N(\gbuff[22][6] ), .A1N(n1542), 
        .Y(n856) );
  OAI2BB2XL U1368 ( .B0(n1497), .B1(n1540), .A0N(\gbuff[22][7] ), .A1N(n1542), 
        .Y(n857) );
  OAI2BB2XL U1369 ( .B0(n1495), .B1(n1540), .A0N(\gbuff[22][8] ), .A1N(n1542), 
        .Y(n858) );
  OAI2BB2XL U1370 ( .B0(n1493), .B1(n1540), .A0N(\gbuff[22][9] ), .A1N(n1542), 
        .Y(n859) );
  OAI2BB2XL U1371 ( .B0(n1491), .B1(n1540), .A0N(\gbuff[22][10] ), .A1N(n1542), 
        .Y(n860) );
  OAI2BB2XL U1372 ( .B0(n1489), .B1(n1540), .A0N(\gbuff[22][11] ), .A1N(n1542), 
        .Y(n861) );
  OAI2BB2XL U1373 ( .B0(n1487), .B1(n1540), .A0N(\gbuff[22][12] ), .A1N(n1542), 
        .Y(n862) );
  OAI2BB2XL U1374 ( .B0(n1485), .B1(n1540), .A0N(\gbuff[22][13] ), .A1N(n1542), 
        .Y(n863) );
  OAI2BB2XL U1375 ( .B0(n1483), .B1(n1541), .A0N(\gbuff[22][14] ), .A1N(n1542), 
        .Y(n864) );
  OAI2BB2XL U1376 ( .B0(n1481), .B1(n1540), .A0N(\gbuff[22][15] ), .A1N(n1541), 
        .Y(n865) );
  OAI2BB2XL U1377 ( .B0(n1479), .B1(n1541), .A0N(\gbuff[22][16] ), .A1N(n1542), 
        .Y(n866) );
  OAI2BB2XL U1378 ( .B0(n1477), .B1(n1540), .A0N(\gbuff[22][17] ), .A1N(n1541), 
        .Y(n867) );
  OAI2BB2XL U1379 ( .B0(n1475), .B1(n1541), .A0N(\gbuff[22][18] ), .A1N(n1541), 
        .Y(n868) );
  OAI2BB2XL U1380 ( .B0(n1473), .B1(n1540), .A0N(\gbuff[22][19] ), .A1N(n1541), 
        .Y(n869) );
  OAI2BB2XL U1381 ( .B0(n1471), .B1(n1541), .A0N(\gbuff[22][20] ), .A1N(n1541), 
        .Y(n870) );
  OAI2BB2XL U1382 ( .B0(n1469), .B1(n1540), .A0N(\gbuff[22][21] ), .A1N(n1541), 
        .Y(n871) );
  OAI2BB2XL U1383 ( .B0(n1467), .B1(n1541), .A0N(\gbuff[22][22] ), .A1N(n1542), 
        .Y(n872) );
  OAI2BB2XL U1384 ( .B0(n1465), .B1(n1541), .A0N(\gbuff[22][23] ), .A1N(n1541), 
        .Y(n873) );
  OAI2BB2XL U1385 ( .B0(n1463), .B1(n135), .A0N(\gbuff[22][24] ), .A1N(n1542), 
        .Y(n874) );
  OAI2BB2XL U1386 ( .B0(n1461), .B1(n1541), .A0N(\gbuff[22][25] ), .A1N(n1542), 
        .Y(n875) );
  OAI2BB2XL U1387 ( .B0(n1459), .B1(n1541), .A0N(\gbuff[22][26] ), .A1N(n1542), 
        .Y(n876) );
  OAI2BB2XL U1388 ( .B0(n1457), .B1(n1541), .A0N(\gbuff[22][27] ), .A1N(n1542), 
        .Y(n877) );
  OAI2BB2XL U1389 ( .B0(n1455), .B1(n1541), .A0N(\gbuff[22][28] ), .A1N(n1542), 
        .Y(n878) );
  OAI2BB2XL U1390 ( .B0(n1453), .B1(n1541), .A0N(\gbuff[22][29] ), .A1N(n1542), 
        .Y(n879) );
  OAI2BB2XL U1391 ( .B0(n1451), .B1(n1541), .A0N(\gbuff[22][30] ), .A1N(n1542), 
        .Y(n880) );
  OAI2BB2XL U1392 ( .B0(n1449), .B1(n1541), .A0N(\gbuff[22][31] ), .A1N(n1540), 
        .Y(n881) );
  OAI2BB2XL U1393 ( .B0(n1511), .B1(n1537), .A0N(\gbuff[23][0] ), .A1N(n1539), 
        .Y(n882) );
  OAI2BB2XL U1394 ( .B0(n1509), .B1(n1537), .A0N(\gbuff[23][1] ), .A1N(n136), 
        .Y(n883) );
  OAI2BB2XL U1395 ( .B0(n1507), .B1(n1537), .A0N(\gbuff[23][2] ), .A1N(n1537), 
        .Y(n884) );
  OAI2BB2XL U1396 ( .B0(n1505), .B1(n1537), .A0N(\gbuff[23][3] ), .A1N(n1539), 
        .Y(n885) );
  OAI2BB2XL U1397 ( .B0(n1503), .B1(n1537), .A0N(\gbuff[23][4] ), .A1N(n1539), 
        .Y(n886) );
  OAI2BB2XL U1398 ( .B0(n1501), .B1(n1537), .A0N(\gbuff[23][5] ), .A1N(n1539), 
        .Y(n887) );
  OAI2BB2XL U1399 ( .B0(n1499), .B1(n1537), .A0N(\gbuff[23][6] ), .A1N(n1539), 
        .Y(n888) );
  OAI2BB2XL U1400 ( .B0(n1497), .B1(n1537), .A0N(\gbuff[23][7] ), .A1N(n1539), 
        .Y(n889) );
  OAI2BB2XL U1401 ( .B0(n1495), .B1(n1537), .A0N(\gbuff[23][8] ), .A1N(n1539), 
        .Y(n890) );
  OAI2BB2XL U1402 ( .B0(n1493), .B1(n1537), .A0N(\gbuff[23][9] ), .A1N(n1539), 
        .Y(n891) );
  OAI2BB2XL U1403 ( .B0(n1491), .B1(n1537), .A0N(\gbuff[23][10] ), .A1N(n1539), 
        .Y(n892) );
  OAI2BB2XL U1404 ( .B0(n1489), .B1(n1537), .A0N(\gbuff[23][11] ), .A1N(n1539), 
        .Y(n893) );
  OAI2BB2XL U1405 ( .B0(n1487), .B1(n1537), .A0N(\gbuff[23][12] ), .A1N(n1539), 
        .Y(n894) );
  OAI2BB2XL U1406 ( .B0(n1485), .B1(n1537), .A0N(\gbuff[23][13] ), .A1N(n1539), 
        .Y(n895) );
  OAI2BB2XL U1407 ( .B0(n1483), .B1(n1538), .A0N(\gbuff[23][14] ), .A1N(n1539), 
        .Y(n896) );
  OAI2BB2XL U1408 ( .B0(n1481), .B1(n1537), .A0N(\gbuff[23][15] ), .A1N(n1538), 
        .Y(n897) );
  OAI2BB2XL U1409 ( .B0(n1479), .B1(n1538), .A0N(\gbuff[23][16] ), .A1N(n1539), 
        .Y(n898) );
  OAI2BB2XL U1410 ( .B0(n1477), .B1(n1537), .A0N(\gbuff[23][17] ), .A1N(n1538), 
        .Y(n899) );
  OAI2BB2XL U1411 ( .B0(n1475), .B1(n1538), .A0N(\gbuff[23][18] ), .A1N(n1538), 
        .Y(n900) );
  OAI2BB2XL U1412 ( .B0(n1473), .B1(n1537), .A0N(\gbuff[23][19] ), .A1N(n1538), 
        .Y(n901) );
  OAI2BB2XL U1413 ( .B0(n1471), .B1(n1538), .A0N(\gbuff[23][20] ), .A1N(n1538), 
        .Y(n902) );
  OAI2BB2XL U1414 ( .B0(n1469), .B1(n1537), .A0N(\gbuff[23][21] ), .A1N(n1538), 
        .Y(n903) );
  OAI2BB2XL U1415 ( .B0(n1467), .B1(n1538), .A0N(\gbuff[23][22] ), .A1N(n1539), 
        .Y(n904) );
  OAI2BB2XL U1416 ( .B0(n1465), .B1(n1538), .A0N(\gbuff[23][23] ), .A1N(n1538), 
        .Y(n905) );
  OAI2BB2XL U1417 ( .B0(n1463), .B1(n136), .A0N(\gbuff[23][24] ), .A1N(n1539), 
        .Y(n906) );
  OAI2BB2XL U1418 ( .B0(n1461), .B1(n1538), .A0N(\gbuff[23][25] ), .A1N(n1539), 
        .Y(n907) );
  OAI2BB2XL U1419 ( .B0(n1459), .B1(n1538), .A0N(\gbuff[23][26] ), .A1N(n1539), 
        .Y(n908) );
  OAI2BB2XL U1420 ( .B0(n1457), .B1(n1538), .A0N(\gbuff[23][27] ), .A1N(n1539), 
        .Y(n909) );
  OAI2BB2XL U1421 ( .B0(n1455), .B1(n1538), .A0N(\gbuff[23][28] ), .A1N(n1539), 
        .Y(n910) );
  OAI2BB2XL U1422 ( .B0(n1453), .B1(n1538), .A0N(\gbuff[23][29] ), .A1N(n1539), 
        .Y(n911) );
  OAI2BB2XL U1423 ( .B0(n1451), .B1(n1538), .A0N(\gbuff[23][30] ), .A1N(n1539), 
        .Y(n912) );
  OAI2BB2XL U1424 ( .B0(n1449), .B1(n1538), .A0N(\gbuff[23][31] ), .A1N(n1537), 
        .Y(n913) );
  OAI2BB2XL U1425 ( .B0(n1511), .B1(n1534), .A0N(\gbuff[24][0] ), .A1N(n1536), 
        .Y(n914) );
  OAI2BB2XL U1426 ( .B0(n1509), .B1(n1534), .A0N(\gbuff[24][1] ), .A1N(n1535), 
        .Y(n915) );
  OAI2BB2XL U1427 ( .B0(n1507), .B1(n1534), .A0N(\gbuff[24][2] ), .A1N(n1534), 
        .Y(n916) );
  OAI2BB2XL U1428 ( .B0(n1505), .B1(n1534), .A0N(\gbuff[24][3] ), .A1N(n1536), 
        .Y(n917) );
  OAI2BB2XL U1429 ( .B0(n1503), .B1(n1534), .A0N(\gbuff[24][4] ), .A1N(n1536), 
        .Y(n918) );
  OAI2BB2XL U1430 ( .B0(n1501), .B1(n1534), .A0N(\gbuff[24][5] ), .A1N(n1536), 
        .Y(n919) );
  OAI2BB2XL U1431 ( .B0(n1499), .B1(n1534), .A0N(\gbuff[24][6] ), .A1N(n1536), 
        .Y(n920) );
  OAI2BB2XL U1432 ( .B0(n1497), .B1(n1534), .A0N(\gbuff[24][7] ), .A1N(n1536), 
        .Y(n921) );
  OAI2BB2XL U1433 ( .B0(n1495), .B1(n1534), .A0N(\gbuff[24][8] ), .A1N(n1536), 
        .Y(n922) );
  OAI2BB2XL U1434 ( .B0(n1493), .B1(n1534), .A0N(\gbuff[24][9] ), .A1N(n1536), 
        .Y(n923) );
  OAI2BB2XL U1435 ( .B0(n1491), .B1(n1534), .A0N(\gbuff[24][10] ), .A1N(n1536), 
        .Y(n924) );
  OAI2BB2XL U1436 ( .B0(n1489), .B1(n1534), .A0N(\gbuff[24][11] ), .A1N(n1536), 
        .Y(n925) );
  OAI2BB2XL U1437 ( .B0(n1487), .B1(n1534), .A0N(\gbuff[24][12] ), .A1N(n1536), 
        .Y(n926) );
  OAI2BB2XL U1438 ( .B0(n1485), .B1(n1534), .A0N(\gbuff[24][13] ), .A1N(n1536), 
        .Y(n927) );
  OAI2BB2XL U1439 ( .B0(n1483), .B1(n1535), .A0N(\gbuff[24][14] ), .A1N(n1536), 
        .Y(n928) );
  OAI2BB2XL U1440 ( .B0(n1481), .B1(n1534), .A0N(\gbuff[24][15] ), .A1N(n1535), 
        .Y(n929) );
  OAI2BB2XL U1441 ( .B0(n1479), .B1(n1535), .A0N(\gbuff[24][16] ), .A1N(n1536), 
        .Y(n930) );
  OAI2BB2XL U1442 ( .B0(n1477), .B1(n1534), .A0N(\gbuff[24][17] ), .A1N(n1535), 
        .Y(n931) );
  OAI2BB2XL U1443 ( .B0(n1475), .B1(n1535), .A0N(\gbuff[24][18] ), .A1N(n1535), 
        .Y(n932) );
  OAI2BB2XL U1444 ( .B0(n1473), .B1(n1534), .A0N(\gbuff[24][19] ), .A1N(n1535), 
        .Y(n933) );
  OAI2BB2XL U1445 ( .B0(n1471), .B1(n1535), .A0N(\gbuff[24][20] ), .A1N(n1535), 
        .Y(n934) );
  OAI2BB2XL U1446 ( .B0(n1469), .B1(n1534), .A0N(\gbuff[24][21] ), .A1N(n1535), 
        .Y(n935) );
  OAI2BB2XL U1447 ( .B0(n1467), .B1(n1535), .A0N(\gbuff[24][22] ), .A1N(n1536), 
        .Y(n936) );
  OAI2BB2XL U1448 ( .B0(n1465), .B1(n1535), .A0N(\gbuff[24][23] ), .A1N(n1535), 
        .Y(n937) );
  OAI2BB2XL U1449 ( .B0(n1463), .B1(n1534), .A0N(\gbuff[24][24] ), .A1N(n1536), 
        .Y(n938) );
  OAI2BB2XL U1450 ( .B0(n1461), .B1(n1535), .A0N(\gbuff[24][25] ), .A1N(n1536), 
        .Y(n939) );
  OAI2BB2XL U1451 ( .B0(n1459), .B1(n1535), .A0N(\gbuff[24][26] ), .A1N(n1536), 
        .Y(n940) );
  OAI2BB2XL U1452 ( .B0(n1457), .B1(n1535), .A0N(\gbuff[24][27] ), .A1N(n1536), 
        .Y(n941) );
  OAI2BB2XL U1453 ( .B0(n1455), .B1(n1535), .A0N(\gbuff[24][28] ), .A1N(n1536), 
        .Y(n942) );
  OAI2BB2XL U1454 ( .B0(n1453), .B1(n1535), .A0N(\gbuff[24][29] ), .A1N(n1536), 
        .Y(n943) );
  OAI2BB2XL U1455 ( .B0(n1451), .B1(n1535), .A0N(\gbuff[24][30] ), .A1N(n1536), 
        .Y(n944) );
  OAI2BB2XL U1456 ( .B0(n1449), .B1(n1535), .A0N(\gbuff[24][31] ), .A1N(n1534), 
        .Y(n945) );
  OAI2BB2XL U1457 ( .B0(n1511), .B1(n1531), .A0N(\gbuff[25][0] ), .A1N(n1533), 
        .Y(n946) );
  OAI2BB2XL U1458 ( .B0(n1509), .B1(n1531), .A0N(\gbuff[25][1] ), .A1N(n1532), 
        .Y(n947) );
  OAI2BB2XL U1459 ( .B0(n1507), .B1(n1531), .A0N(\gbuff[25][2] ), .A1N(n1531), 
        .Y(n948) );
  OAI2BB2XL U1460 ( .B0(n1505), .B1(n1531), .A0N(\gbuff[25][3] ), .A1N(n1533), 
        .Y(n949) );
  OAI2BB2XL U1461 ( .B0(n1503), .B1(n1531), .A0N(\gbuff[25][4] ), .A1N(n1533), 
        .Y(n950) );
  OAI2BB2XL U1462 ( .B0(n1501), .B1(n1531), .A0N(\gbuff[25][5] ), .A1N(n1533), 
        .Y(n951) );
  OAI2BB2XL U1463 ( .B0(n1499), .B1(n1531), .A0N(\gbuff[25][6] ), .A1N(n1533), 
        .Y(n952) );
  OAI2BB2XL U1464 ( .B0(n1497), .B1(n1531), .A0N(\gbuff[25][7] ), .A1N(n1533), 
        .Y(n953) );
  OAI2BB2XL U1465 ( .B0(n1495), .B1(n1531), .A0N(\gbuff[25][8] ), .A1N(n1533), 
        .Y(n954) );
  OAI2BB2XL U1466 ( .B0(n1493), .B1(n1531), .A0N(\gbuff[25][9] ), .A1N(n1533), 
        .Y(n955) );
  OAI2BB2XL U1467 ( .B0(n1491), .B1(n1531), .A0N(\gbuff[25][10] ), .A1N(n1533), 
        .Y(n956) );
  OAI2BB2XL U1468 ( .B0(n1489), .B1(n1531), .A0N(\gbuff[25][11] ), .A1N(n1533), 
        .Y(n957) );
  OAI2BB2XL U1469 ( .B0(n1487), .B1(n1531), .A0N(\gbuff[25][12] ), .A1N(n1533), 
        .Y(n958) );
  OAI2BB2XL U1470 ( .B0(n1485), .B1(n1531), .A0N(\gbuff[25][13] ), .A1N(n1533), 
        .Y(n959) );
  OAI2BB2XL U1471 ( .B0(n1483), .B1(n1532), .A0N(\gbuff[25][14] ), .A1N(n1533), 
        .Y(n960) );
  OAI2BB2XL U1472 ( .B0(n1481), .B1(n1531), .A0N(\gbuff[25][15] ), .A1N(n1532), 
        .Y(n961) );
  OAI2BB2XL U1473 ( .B0(n1479), .B1(n1532), .A0N(\gbuff[25][16] ), .A1N(n1533), 
        .Y(n962) );
  OAI2BB2XL U1474 ( .B0(n1477), .B1(n1531), .A0N(\gbuff[25][17] ), .A1N(n1532), 
        .Y(n963) );
  OAI2BB2XL U1475 ( .B0(n1475), .B1(n1532), .A0N(\gbuff[25][18] ), .A1N(n1532), 
        .Y(n964) );
  OAI2BB2XL U1476 ( .B0(n1473), .B1(n1531), .A0N(\gbuff[25][19] ), .A1N(n1532), 
        .Y(n965) );
  OAI2BB2XL U1477 ( .B0(n1471), .B1(n1532), .A0N(\gbuff[25][20] ), .A1N(n1532), 
        .Y(n966) );
  OAI2BB2XL U1478 ( .B0(n1469), .B1(n1531), .A0N(\gbuff[25][21] ), .A1N(n1532), 
        .Y(n967) );
  OAI2BB2XL U1479 ( .B0(n1467), .B1(n1532), .A0N(\gbuff[25][22] ), .A1N(n1533), 
        .Y(n968) );
  OAI2BB2XL U1480 ( .B0(n1465), .B1(n1532), .A0N(\gbuff[25][23] ), .A1N(n1532), 
        .Y(n969) );
  OAI2BB2XL U1481 ( .B0(n1463), .B1(n1531), .A0N(\gbuff[25][24] ), .A1N(n1533), 
        .Y(n970) );
  OAI2BB2XL U1482 ( .B0(n1461), .B1(n1532), .A0N(\gbuff[25][25] ), .A1N(n1533), 
        .Y(n971) );
  OAI2BB2XL U1483 ( .B0(n1459), .B1(n1532), .A0N(\gbuff[25][26] ), .A1N(n1533), 
        .Y(n972) );
  OAI2BB2XL U1484 ( .B0(n1457), .B1(n1532), .A0N(\gbuff[25][27] ), .A1N(n1533), 
        .Y(n973) );
  OAI2BB2XL U1485 ( .B0(n1455), .B1(n1532), .A0N(\gbuff[25][28] ), .A1N(n1533), 
        .Y(n974) );
  OAI2BB2XL U1486 ( .B0(n1453), .B1(n1532), .A0N(\gbuff[25][29] ), .A1N(n1533), 
        .Y(n975) );
  OAI2BB2XL U1487 ( .B0(n1451), .B1(n1532), .A0N(\gbuff[25][30] ), .A1N(n1533), 
        .Y(n976) );
  OAI2BB2XL U1488 ( .B0(n1449), .B1(n1532), .A0N(\gbuff[25][31] ), .A1N(n1531), 
        .Y(n977) );
  OAI2BB2XL U1489 ( .B0(n1511), .B1(n1528), .A0N(\gbuff[26][0] ), .A1N(n1530), 
        .Y(n978) );
  OAI2BB2XL U1490 ( .B0(n1509), .B1(n1528), .A0N(\gbuff[26][1] ), .A1N(n1529), 
        .Y(n979) );
  OAI2BB2XL U1491 ( .B0(n1507), .B1(n1528), .A0N(\gbuff[26][2] ), .A1N(n1528), 
        .Y(n980) );
  OAI2BB2XL U1492 ( .B0(n1505), .B1(n1528), .A0N(\gbuff[26][3] ), .A1N(n1530), 
        .Y(n981) );
  OAI2BB2XL U1493 ( .B0(n1503), .B1(n1528), .A0N(\gbuff[26][4] ), .A1N(n1530), 
        .Y(n982) );
  OAI2BB2XL U1494 ( .B0(n1501), .B1(n1528), .A0N(\gbuff[26][5] ), .A1N(n1530), 
        .Y(n983) );
  OAI2BB2XL U1495 ( .B0(n1499), .B1(n1528), .A0N(\gbuff[26][6] ), .A1N(n1530), 
        .Y(n984) );
  OAI2BB2XL U1496 ( .B0(n1497), .B1(n1528), .A0N(\gbuff[26][7] ), .A1N(n1530), 
        .Y(n985) );
  OAI2BB2XL U1497 ( .B0(n1495), .B1(n1528), .A0N(\gbuff[26][8] ), .A1N(n1530), 
        .Y(n986) );
  OAI2BB2XL U1498 ( .B0(n1493), .B1(n1528), .A0N(\gbuff[26][9] ), .A1N(n1530), 
        .Y(n987) );
  OAI2BB2XL U1499 ( .B0(n1491), .B1(n1528), .A0N(\gbuff[26][10] ), .A1N(n1530), 
        .Y(n988) );
  OAI2BB2XL U1500 ( .B0(n1489), .B1(n1528), .A0N(\gbuff[26][11] ), .A1N(n1530), 
        .Y(n989) );
  OAI2BB2XL U1501 ( .B0(n1487), .B1(n1528), .A0N(\gbuff[26][12] ), .A1N(n1530), 
        .Y(n990) );
  OAI2BB2XL U1502 ( .B0(n1485), .B1(n1528), .A0N(\gbuff[26][13] ), .A1N(n1530), 
        .Y(n991) );
  OAI2BB2XL U1503 ( .B0(n1483), .B1(n1529), .A0N(\gbuff[26][14] ), .A1N(n1530), 
        .Y(n992) );
  OAI2BB2XL U1504 ( .B0(n1481), .B1(n1528), .A0N(\gbuff[26][15] ), .A1N(n1529), 
        .Y(n993) );
  OAI2BB2XL U1505 ( .B0(n1479), .B1(n1529), .A0N(\gbuff[26][16] ), .A1N(n1530), 
        .Y(n994) );
  OAI2BB2XL U1506 ( .B0(n1477), .B1(n1528), .A0N(\gbuff[26][17] ), .A1N(n1529), 
        .Y(n995) );
  OAI2BB2XL U1507 ( .B0(n1475), .B1(n1529), .A0N(\gbuff[26][18] ), .A1N(n1529), 
        .Y(n996) );
  OAI2BB2XL U1508 ( .B0(n1473), .B1(n1528), .A0N(\gbuff[26][19] ), .A1N(n1529), 
        .Y(n997) );
  OAI2BB2XL U1509 ( .B0(n1471), .B1(n1529), .A0N(\gbuff[26][20] ), .A1N(n1529), 
        .Y(n998) );
  OAI2BB2XL U1510 ( .B0(n1469), .B1(n1528), .A0N(\gbuff[26][21] ), .A1N(n1529), 
        .Y(n999) );
  OAI2BB2XL U1511 ( .B0(n1467), .B1(n1529), .A0N(\gbuff[26][22] ), .A1N(n1530), 
        .Y(n1000) );
  OAI2BB2XL U1512 ( .B0(n1465), .B1(n1529), .A0N(\gbuff[26][23] ), .A1N(n1529), 
        .Y(n1001) );
  OAI2BB2XL U1513 ( .B0(n1463), .B1(n1528), .A0N(\gbuff[26][24] ), .A1N(n1530), 
        .Y(n1002) );
  OAI2BB2XL U1514 ( .B0(n1461), .B1(n1529), .A0N(\gbuff[26][25] ), .A1N(n1530), 
        .Y(n1003) );
  OAI2BB2XL U1515 ( .B0(n1459), .B1(n1529), .A0N(\gbuff[26][26] ), .A1N(n1530), 
        .Y(n1004) );
  OAI2BB2XL U1516 ( .B0(n1457), .B1(n1529), .A0N(\gbuff[26][27] ), .A1N(n1530), 
        .Y(n1005) );
  OAI2BB2XL U1517 ( .B0(n1455), .B1(n1529), .A0N(\gbuff[26][28] ), .A1N(n1530), 
        .Y(n1006) );
  OAI2BB2XL U1518 ( .B0(n1453), .B1(n1529), .A0N(\gbuff[26][29] ), .A1N(n1530), 
        .Y(n1007) );
  OAI2BB2XL U1519 ( .B0(n1451), .B1(n1529), .A0N(\gbuff[26][30] ), .A1N(n1530), 
        .Y(n1008) );
  OAI2BB2XL U1520 ( .B0(n1449), .B1(n1529), .A0N(\gbuff[26][31] ), .A1N(n1528), 
        .Y(n1009) );
  OAI2BB2XL U1521 ( .B0(n1511), .B1(n1525), .A0N(\gbuff[27][0] ), .A1N(n1527), 
        .Y(n1010) );
  OAI2BB2XL U1522 ( .B0(n1509), .B1(n1525), .A0N(\gbuff[27][1] ), .A1N(n1526), 
        .Y(n1011) );
  OAI2BB2XL U1523 ( .B0(n1507), .B1(n1525), .A0N(\gbuff[27][2] ), .A1N(n1525), 
        .Y(n1012) );
  OAI2BB2XL U1524 ( .B0(n1505), .B1(n1525), .A0N(\gbuff[27][3] ), .A1N(n1527), 
        .Y(n1013) );
  OAI2BB2XL U1525 ( .B0(n1503), .B1(n1525), .A0N(\gbuff[27][4] ), .A1N(n1527), 
        .Y(n1014) );
  OAI2BB2XL U1526 ( .B0(n1501), .B1(n1525), .A0N(\gbuff[27][5] ), .A1N(n1527), 
        .Y(n1015) );
  OAI2BB2XL U1527 ( .B0(n1499), .B1(n1525), .A0N(\gbuff[27][6] ), .A1N(n1527), 
        .Y(n1016) );
  OAI2BB2XL U1528 ( .B0(n1497), .B1(n1525), .A0N(\gbuff[27][7] ), .A1N(n1527), 
        .Y(n1017) );
  OAI2BB2XL U1529 ( .B0(n1495), .B1(n1525), .A0N(\gbuff[27][8] ), .A1N(n1527), 
        .Y(n1018) );
  OAI2BB2XL U1530 ( .B0(n1493), .B1(n1525), .A0N(\gbuff[27][9] ), .A1N(n1527), 
        .Y(n1019) );
  OAI2BB2XL U1531 ( .B0(n1491), .B1(n1525), .A0N(\gbuff[27][10] ), .A1N(n1527), 
        .Y(n1020) );
  OAI2BB2XL U1532 ( .B0(n1489), .B1(n1525), .A0N(\gbuff[27][11] ), .A1N(n1527), 
        .Y(n1021) );
  OAI2BB2XL U1533 ( .B0(n1487), .B1(n1525), .A0N(\gbuff[27][12] ), .A1N(n1527), 
        .Y(n1022) );
  OAI2BB2XL U1534 ( .B0(n1485), .B1(n1525), .A0N(\gbuff[27][13] ), .A1N(n1527), 
        .Y(n1023) );
  OAI2BB2XL U1535 ( .B0(n1483), .B1(n1526), .A0N(\gbuff[27][14] ), .A1N(n1527), 
        .Y(n1024) );
  OAI2BB2XL U1536 ( .B0(n1481), .B1(n1525), .A0N(\gbuff[27][15] ), .A1N(n1526), 
        .Y(n1025) );
  OAI2BB2XL U1537 ( .B0(n1479), .B1(n1526), .A0N(\gbuff[27][16] ), .A1N(n1527), 
        .Y(n1026) );
  OAI2BB2XL U1538 ( .B0(n1477), .B1(n1525), .A0N(\gbuff[27][17] ), .A1N(n1526), 
        .Y(n1027) );
  OAI2BB2XL U1539 ( .B0(n1475), .B1(n1526), .A0N(\gbuff[27][18] ), .A1N(n1526), 
        .Y(n1028) );
  OAI2BB2XL U1540 ( .B0(n1473), .B1(n1525), .A0N(\gbuff[27][19] ), .A1N(n1526), 
        .Y(n1029) );
  OAI2BB2XL U1541 ( .B0(n1471), .B1(n1526), .A0N(\gbuff[27][20] ), .A1N(n1526), 
        .Y(n1030) );
  OAI2BB2XL U1542 ( .B0(n1469), .B1(n1525), .A0N(\gbuff[27][21] ), .A1N(n1526), 
        .Y(n1031) );
  OAI2BB2XL U1543 ( .B0(n1467), .B1(n1526), .A0N(\gbuff[27][22] ), .A1N(n1527), 
        .Y(n1032) );
  OAI2BB2XL U1544 ( .B0(n1465), .B1(n1526), .A0N(\gbuff[27][23] ), .A1N(n1526), 
        .Y(n1033) );
  OAI2BB2XL U1545 ( .B0(n1463), .B1(n1525), .A0N(\gbuff[27][24] ), .A1N(n1527), 
        .Y(n1034) );
  OAI2BB2XL U1546 ( .B0(n1461), .B1(n1526), .A0N(\gbuff[27][25] ), .A1N(n1527), 
        .Y(n1035) );
  OAI2BB2XL U1547 ( .B0(n1459), .B1(n1526), .A0N(\gbuff[27][26] ), .A1N(n1527), 
        .Y(n1036) );
  OAI2BB2XL U1548 ( .B0(n1457), .B1(n1526), .A0N(\gbuff[27][27] ), .A1N(n1527), 
        .Y(n1037) );
  OAI2BB2XL U1549 ( .B0(n1455), .B1(n1526), .A0N(\gbuff[27][28] ), .A1N(n1527), 
        .Y(n1038) );
  OAI2BB2XL U1550 ( .B0(n1453), .B1(n1526), .A0N(\gbuff[27][29] ), .A1N(n1527), 
        .Y(n1039) );
  OAI2BB2XL U1551 ( .B0(n1451), .B1(n1526), .A0N(\gbuff[27][30] ), .A1N(n1527), 
        .Y(n1040) );
  OAI2BB2XL U1552 ( .B0(n1449), .B1(n1526), .A0N(\gbuff[27][31] ), .A1N(n1525), 
        .Y(n1041) );
  OAI2BB2XL U1553 ( .B0(n1511), .B1(n1523), .A0N(\gbuff[28][0] ), .A1N(n1523), 
        .Y(n1042) );
  OAI2BB2XL U1554 ( .B0(n1509), .B1(n1522), .A0N(\gbuff[28][1] ), .A1N(n1522), 
        .Y(n1043) );
  OAI2BB2XL U1555 ( .B0(n1507), .B1(n1522), .A0N(\gbuff[28][2] ), .A1N(n1523), 
        .Y(n1044) );
  OAI2BB2XL U1556 ( .B0(n1505), .B1(n1522), .A0N(\gbuff[28][3] ), .A1N(n1524), 
        .Y(n1045) );
  OAI2BB2XL U1557 ( .B0(n1503), .B1(n1522), .A0N(\gbuff[28][4] ), .A1N(n1522), 
        .Y(n1046) );
  OAI2BB2XL U1558 ( .B0(n1501), .B1(n1522), .A0N(\gbuff[28][5] ), .A1N(n1524), 
        .Y(n1047) );
  OAI2BB2XL U1559 ( .B0(n1499), .B1(n1522), .A0N(\gbuff[28][6] ), .A1N(n1524), 
        .Y(n1048) );
  OAI2BB2XL U1560 ( .B0(n1497), .B1(n1522), .A0N(\gbuff[28][7] ), .A1N(n1524), 
        .Y(n1049) );
  OAI2BB2XL U1561 ( .B0(n1495), .B1(n1522), .A0N(\gbuff[28][8] ), .A1N(n1524), 
        .Y(n1050) );
  OAI2BB2XL U1562 ( .B0(n1493), .B1(n1522), .A0N(\gbuff[28][9] ), .A1N(n1524), 
        .Y(n1051) );
  OAI2BB2XL U1563 ( .B0(n1491), .B1(n1522), .A0N(\gbuff[28][10] ), .A1N(n1524), 
        .Y(n1052) );
  OAI2BB2XL U1564 ( .B0(n1489), .B1(n1522), .A0N(\gbuff[28][11] ), .A1N(n1524), 
        .Y(n1053) );
  OAI2BB2XL U1565 ( .B0(n1487), .B1(n1522), .A0N(\gbuff[28][12] ), .A1N(n1524), 
        .Y(n1054) );
  OAI2BB2XL U1566 ( .B0(n1485), .B1(n1523), .A0N(\gbuff[28][13] ), .A1N(n1524), 
        .Y(n1055) );
  OAI2BB2XL U1567 ( .B0(n1483), .B1(n1523), .A0N(\gbuff[28][14] ), .A1N(n1524), 
        .Y(n1056) );
  OAI2BB2XL U1568 ( .B0(n1481), .B1(n1523), .A0N(\gbuff[28][15] ), .A1N(n1524), 
        .Y(n1057) );
  OAI2BB2XL U1569 ( .B0(n1479), .B1(n1523), .A0N(\gbuff[28][16] ), .A1N(n1524), 
        .Y(n1058) );
  OAI2BB2XL U1570 ( .B0(n1477), .B1(n1523), .A0N(\gbuff[28][17] ), .A1N(n1524), 
        .Y(n1059) );
  OAI2BB2XL U1571 ( .B0(n1475), .B1(n1523), .A0N(\gbuff[28][18] ), .A1N(n142), 
        .Y(n1060) );
  OAI2BB2XL U1572 ( .B0(n1473), .B1(n1523), .A0N(\gbuff[28][19] ), .A1N(n1522), 
        .Y(n1061) );
  OAI2BB2XL U1573 ( .B0(n1471), .B1(n1523), .A0N(\gbuff[28][20] ), .A1N(n1523), 
        .Y(n1062) );
  OAI2BB2XL U1574 ( .B0(n1469), .B1(n1523), .A0N(\gbuff[28][21] ), .A1N(n142), 
        .Y(n1063) );
  OAI2BB2XL U1575 ( .B0(n1467), .B1(n1523), .A0N(\gbuff[28][22] ), .A1N(n1524), 
        .Y(n1064) );
  OAI2BB2XL U1576 ( .B0(n1465), .B1(n1522), .A0N(\gbuff[28][23] ), .A1N(n1524), 
        .Y(n1065) );
  OAI2BB2XL U1577 ( .B0(n1463), .B1(n1523), .A0N(\gbuff[28][24] ), .A1N(n1524), 
        .Y(n1066) );
  OAI2BB2XL U1578 ( .B0(n1461), .B1(n1523), .A0N(\gbuff[28][25] ), .A1N(n1524), 
        .Y(n1067) );
  OAI2BB2XL U1579 ( .B0(n1459), .B1(n1522), .A0N(\gbuff[28][26] ), .A1N(n1524), 
        .Y(n1068) );
  OAI2BB2XL U1580 ( .B0(n1457), .B1(n1523), .A0N(\gbuff[28][27] ), .A1N(n1524), 
        .Y(n1069) );
  OAI2BB2XL U1581 ( .B0(n1455), .B1(n1522), .A0N(\gbuff[28][28] ), .A1N(n1524), 
        .Y(n1070) );
  OAI2BB2XL U1582 ( .B0(n1453), .B1(n1523), .A0N(\gbuff[28][29] ), .A1N(n1524), 
        .Y(n1071) );
  OAI2BB2XL U1583 ( .B0(n1451), .B1(n1522), .A0N(\gbuff[28][30] ), .A1N(n1523), 
        .Y(n1072) );
  OAI2BB2XL U1584 ( .B0(n1449), .B1(n1523), .A0N(\gbuff[28][31] ), .A1N(n1522), 
        .Y(n1073) );
  OAI2BB2XL U1585 ( .B0(n1511), .B1(n1519), .A0N(\gbuff[29][0] ), .A1N(n1521), 
        .Y(n1074) );
  OAI2BB2XL U1586 ( .B0(n1509), .B1(n1519), .A0N(\gbuff[29][1] ), .A1N(n143), 
        .Y(n1075) );
  OAI2BB2XL U1587 ( .B0(n1507), .B1(n1519), .A0N(\gbuff[29][2] ), .A1N(n1519), 
        .Y(n1076) );
  OAI2BB2XL U1588 ( .B0(n1505), .B1(n1519), .A0N(\gbuff[29][3] ), .A1N(n1521), 
        .Y(n1077) );
  OAI2BB2XL U1589 ( .B0(n1503), .B1(n1519), .A0N(\gbuff[29][4] ), .A1N(n1521), 
        .Y(n1078) );
  OAI2BB2XL U1590 ( .B0(n1501), .B1(n1519), .A0N(\gbuff[29][5] ), .A1N(n1521), 
        .Y(n1079) );
  OAI2BB2XL U1591 ( .B0(n1499), .B1(n1519), .A0N(\gbuff[29][6] ), .A1N(n1521), 
        .Y(n1080) );
  OAI2BB2XL U1592 ( .B0(n1497), .B1(n1519), .A0N(\gbuff[29][7] ), .A1N(n1521), 
        .Y(n1081) );
  OAI2BB2XL U1593 ( .B0(n1495), .B1(n1519), .A0N(\gbuff[29][8] ), .A1N(n1521), 
        .Y(n1082) );
  OAI2BB2XL U1594 ( .B0(n1493), .B1(n1519), .A0N(\gbuff[29][9] ), .A1N(n1521), 
        .Y(n1083) );
  OAI2BB2XL U1595 ( .B0(n1491), .B1(n1519), .A0N(\gbuff[29][10] ), .A1N(n1521), 
        .Y(n1084) );
  OAI2BB2XL U1596 ( .B0(n1489), .B1(n1519), .A0N(\gbuff[29][11] ), .A1N(n1521), 
        .Y(n1085) );
  OAI2BB2XL U1597 ( .B0(n1487), .B1(n1519), .A0N(\gbuff[29][12] ), .A1N(n1521), 
        .Y(n1086) );
  OAI2BB2XL U1598 ( .B0(n1485), .B1(n1519), .A0N(\gbuff[29][13] ), .A1N(n1521), 
        .Y(n1087) );
  OAI2BB2XL U1599 ( .B0(n1483), .B1(n1520), .A0N(\gbuff[29][14] ), .A1N(n1521), 
        .Y(n1088) );
  OAI2BB2XL U1600 ( .B0(n1481), .B1(n1519), .A0N(\gbuff[29][15] ), .A1N(n1520), 
        .Y(n1089) );
  OAI2BB2XL U1601 ( .B0(n1479), .B1(n1520), .A0N(\gbuff[29][16] ), .A1N(n1521), 
        .Y(n1090) );
  OAI2BB2XL U1602 ( .B0(n1477), .B1(n1519), .A0N(\gbuff[29][17] ), .A1N(n1520), 
        .Y(n1091) );
  OAI2BB2XL U1603 ( .B0(n1475), .B1(n1520), .A0N(\gbuff[29][18] ), .A1N(n1520), 
        .Y(n1092) );
  OAI2BB2XL U1604 ( .B0(n1473), .B1(n1519), .A0N(\gbuff[29][19] ), .A1N(n1520), 
        .Y(n1093) );
  OAI2BB2XL U1605 ( .B0(n1471), .B1(n1520), .A0N(\gbuff[29][20] ), .A1N(n1520), 
        .Y(n1094) );
  OAI2BB2XL U1606 ( .B0(n1469), .B1(n1519), .A0N(\gbuff[29][21] ), .A1N(n1520), 
        .Y(n1095) );
  OAI2BB2XL U1607 ( .B0(n1467), .B1(n1520), .A0N(\gbuff[29][22] ), .A1N(n1521), 
        .Y(n1096) );
  OAI2BB2XL U1608 ( .B0(n1465), .B1(n1520), .A0N(\gbuff[29][23] ), .A1N(n1520), 
        .Y(n1097) );
  OAI2BB2XL U1609 ( .B0(n1463), .B1(n143), .A0N(\gbuff[29][24] ), .A1N(n1521), 
        .Y(n1098) );
  OAI2BB2XL U1610 ( .B0(n1461), .B1(n1520), .A0N(\gbuff[29][25] ), .A1N(n1521), 
        .Y(n1099) );
  OAI2BB2XL U1611 ( .B0(n1459), .B1(n1520), .A0N(\gbuff[29][26] ), .A1N(n1521), 
        .Y(n1100) );
  OAI2BB2XL U1612 ( .B0(n1457), .B1(n1520), .A0N(\gbuff[29][27] ), .A1N(n1521), 
        .Y(n1101) );
  OAI2BB2XL U1613 ( .B0(n1455), .B1(n1520), .A0N(\gbuff[29][28] ), .A1N(n1521), 
        .Y(n1102) );
  OAI2BB2XL U1614 ( .B0(n1453), .B1(n1520), .A0N(\gbuff[29][29] ), .A1N(n1521), 
        .Y(n1103) );
  OAI2BB2XL U1615 ( .B0(n1451), .B1(n1520), .A0N(\gbuff[29][30] ), .A1N(n1521), 
        .Y(n1104) );
  OAI2BB2XL U1616 ( .B0(n1449), .B1(n1520), .A0N(\gbuff[29][31] ), .A1N(n1519), 
        .Y(n1105) );
  OAI2BB2XL U1617 ( .B0(n1511), .B1(n1516), .A0N(\gbuff[30][0] ), .A1N(n1518), 
        .Y(n1106) );
  OAI2BB2XL U1618 ( .B0(n1509), .B1(n1516), .A0N(\gbuff[30][1] ), .A1N(n144), 
        .Y(n1107) );
  OAI2BB2XL U1619 ( .B0(n1507), .B1(n1516), .A0N(\gbuff[30][2] ), .A1N(n1516), 
        .Y(n1108) );
  OAI2BB2XL U1620 ( .B0(n1505), .B1(n1516), .A0N(\gbuff[30][3] ), .A1N(n1518), 
        .Y(n1109) );
  OAI2BB2XL U1621 ( .B0(n1503), .B1(n1516), .A0N(\gbuff[30][4] ), .A1N(n1518), 
        .Y(n1110) );
  OAI2BB2XL U1622 ( .B0(n1501), .B1(n1516), .A0N(\gbuff[30][5] ), .A1N(n1518), 
        .Y(n1111) );
  OAI2BB2XL U1623 ( .B0(n1499), .B1(n1516), .A0N(\gbuff[30][6] ), .A1N(n1518), 
        .Y(n1112) );
  OAI2BB2XL U1624 ( .B0(n1497), .B1(n1516), .A0N(\gbuff[30][7] ), .A1N(n1518), 
        .Y(n1113) );
  OAI2BB2XL U1625 ( .B0(n1495), .B1(n1516), .A0N(\gbuff[30][8] ), .A1N(n1518), 
        .Y(n1114) );
  OAI2BB2XL U1626 ( .B0(n1493), .B1(n1516), .A0N(\gbuff[30][9] ), .A1N(n1518), 
        .Y(n1115) );
  OAI2BB2XL U1627 ( .B0(n1491), .B1(n1516), .A0N(\gbuff[30][10] ), .A1N(n1518), 
        .Y(n1116) );
  OAI2BB2XL U1628 ( .B0(n1489), .B1(n1516), .A0N(\gbuff[30][11] ), .A1N(n1518), 
        .Y(n1117) );
  OAI2BB2XL U1629 ( .B0(n1487), .B1(n1516), .A0N(\gbuff[30][12] ), .A1N(n1518), 
        .Y(n1118) );
  OAI2BB2XL U1630 ( .B0(n1485), .B1(n1516), .A0N(\gbuff[30][13] ), .A1N(n1518), 
        .Y(n1119) );
  OAI2BB2XL U1631 ( .B0(n1483), .B1(n1517), .A0N(\gbuff[30][14] ), .A1N(n1518), 
        .Y(n1120) );
  OAI2BB2XL U1632 ( .B0(n1481), .B1(n1516), .A0N(\gbuff[30][15] ), .A1N(n1517), 
        .Y(n1121) );
  OAI2BB2XL U1633 ( .B0(n1479), .B1(n1517), .A0N(\gbuff[30][16] ), .A1N(n1518), 
        .Y(n1122) );
  OAI2BB2XL U1634 ( .B0(n1477), .B1(n1516), .A0N(\gbuff[30][17] ), .A1N(n1517), 
        .Y(n1123) );
  OAI2BB2XL U1635 ( .B0(n1475), .B1(n1517), .A0N(\gbuff[30][18] ), .A1N(n1517), 
        .Y(n1124) );
  OAI2BB2XL U1636 ( .B0(n1473), .B1(n1516), .A0N(\gbuff[30][19] ), .A1N(n1517), 
        .Y(n1125) );
  OAI2BB2XL U1637 ( .B0(n1471), .B1(n1517), .A0N(\gbuff[30][20] ), .A1N(n1517), 
        .Y(n1126) );
  OAI2BB2XL U1638 ( .B0(n1469), .B1(n1516), .A0N(\gbuff[30][21] ), .A1N(n1517), 
        .Y(n1127) );
  OAI2BB2XL U1639 ( .B0(n1467), .B1(n1517), .A0N(\gbuff[30][22] ), .A1N(n1518), 
        .Y(n1128) );
  OAI2BB2XL U1640 ( .B0(n1465), .B1(n1517), .A0N(\gbuff[30][23] ), .A1N(n1517), 
        .Y(n1129) );
  OAI2BB2XL U1641 ( .B0(n1463), .B1(n144), .A0N(\gbuff[30][24] ), .A1N(n1518), 
        .Y(n1130) );
  OAI2BB2XL U1642 ( .B0(n1461), .B1(n1517), .A0N(\gbuff[30][25] ), .A1N(n1518), 
        .Y(n1131) );
  OAI2BB2XL U1643 ( .B0(n1459), .B1(n1517), .A0N(\gbuff[30][26] ), .A1N(n1518), 
        .Y(n1132) );
  OAI2BB2XL U1644 ( .B0(n1457), .B1(n1517), .A0N(\gbuff[30][27] ), .A1N(n1518), 
        .Y(n1133) );
  OAI2BB2XL U1645 ( .B0(n1455), .B1(n1517), .A0N(\gbuff[30][28] ), .A1N(n1518), 
        .Y(n1134) );
  OAI2BB2XL U1646 ( .B0(n1453), .B1(n1517), .A0N(\gbuff[30][29] ), .A1N(n1518), 
        .Y(n1135) );
  OAI2BB2XL U1647 ( .B0(n1451), .B1(n1517), .A0N(\gbuff[30][30] ), .A1N(n1518), 
        .Y(n1136) );
  OAI2BB2XL U1648 ( .B0(n1449), .B1(n1517), .A0N(\gbuff[30][31] ), .A1N(n1516), 
        .Y(n1137) );
  OAI2BB2XL U1649 ( .B0(n1511), .B1(n1513), .A0N(\gbuff[31][0] ), .A1N(n1515), 
        .Y(n1138) );
  OAI2BB2XL U1650 ( .B0(n1509), .B1(n1513), .A0N(\gbuff[31][1] ), .A1N(n145), 
        .Y(n1139) );
  OAI2BB2XL U1651 ( .B0(n1507), .B1(n1513), .A0N(\gbuff[31][2] ), .A1N(n1513), 
        .Y(n1140) );
  OAI2BB2XL U1652 ( .B0(n1505), .B1(n1513), .A0N(\gbuff[31][3] ), .A1N(n1515), 
        .Y(n1141) );
  OAI2BB2XL U1653 ( .B0(n1503), .B1(n1513), .A0N(\gbuff[31][4] ), .A1N(n1515), 
        .Y(n1142) );
  OAI2BB2XL U1654 ( .B0(n1501), .B1(n1513), .A0N(\gbuff[31][5] ), .A1N(n1515), 
        .Y(n1143) );
  OAI2BB2XL U1655 ( .B0(n1499), .B1(n1513), .A0N(\gbuff[31][6] ), .A1N(n1515), 
        .Y(n1144) );
  OAI2BB2XL U1656 ( .B0(n1497), .B1(n1513), .A0N(\gbuff[31][7] ), .A1N(n1515), 
        .Y(n1145) );
  OAI2BB2XL U1657 ( .B0(n1495), .B1(n1513), .A0N(\gbuff[31][8] ), .A1N(n1515), 
        .Y(n1146) );
  OAI2BB2XL U1658 ( .B0(n1493), .B1(n1513), .A0N(\gbuff[31][9] ), .A1N(n1515), 
        .Y(n1147) );
  OAI2BB2XL U1659 ( .B0(n1491), .B1(n1513), .A0N(\gbuff[31][10] ), .A1N(n1515), 
        .Y(n1148) );
  OAI2BB2XL U1660 ( .B0(n1489), .B1(n1513), .A0N(\gbuff[31][11] ), .A1N(n1515), 
        .Y(n1149) );
  OAI2BB2XL U1661 ( .B0(n1487), .B1(n1513), .A0N(\gbuff[31][12] ), .A1N(n1515), 
        .Y(n1150) );
  OAI2BB2XL U1662 ( .B0(n1485), .B1(n1513), .A0N(\gbuff[31][13] ), .A1N(n1515), 
        .Y(n1151) );
  OAI2BB2XL U1663 ( .B0(n1483), .B1(n1514), .A0N(\gbuff[31][14] ), .A1N(n1515), 
        .Y(n1152) );
  OAI2BB2XL U1664 ( .B0(n1481), .B1(n1513), .A0N(\gbuff[31][15] ), .A1N(n1514), 
        .Y(n1153) );
  OAI2BB2XL U1665 ( .B0(n1479), .B1(n1514), .A0N(\gbuff[31][16] ), .A1N(n1515), 
        .Y(n1154) );
  OAI2BB2XL U1666 ( .B0(n1477), .B1(n1513), .A0N(\gbuff[31][17] ), .A1N(n1514), 
        .Y(n1155) );
  OAI2BB2XL U1667 ( .B0(n1475), .B1(n1514), .A0N(\gbuff[31][18] ), .A1N(n1514), 
        .Y(n1156) );
  OAI2BB2XL U1668 ( .B0(n1473), .B1(n1513), .A0N(\gbuff[31][19] ), .A1N(n1514), 
        .Y(n1157) );
  OAI2BB2XL U1669 ( .B0(n1471), .B1(n1514), .A0N(\gbuff[31][20] ), .A1N(n1514), 
        .Y(n1158) );
  OAI2BB2XL U1670 ( .B0(n1469), .B1(n1513), .A0N(\gbuff[31][21] ), .A1N(n1514), 
        .Y(n1159) );
  OAI2BB2XL U1671 ( .B0(n1467), .B1(n1514), .A0N(\gbuff[31][22] ), .A1N(n1515), 
        .Y(n1160) );
  OAI2BB2XL U1672 ( .B0(n1465), .B1(n1514), .A0N(\gbuff[31][23] ), .A1N(n1514), 
        .Y(n1161) );
  OAI2BB2XL U1673 ( .B0(n1463), .B1(n145), .A0N(\gbuff[31][24] ), .A1N(n1515), 
        .Y(n1162) );
  OAI2BB2XL U1674 ( .B0(n1461), .B1(n1514), .A0N(\gbuff[31][25] ), .A1N(n1515), 
        .Y(n1163) );
  OAI2BB2XL U1675 ( .B0(n1459), .B1(n1514), .A0N(\gbuff[31][26] ), .A1N(n1515), 
        .Y(n1164) );
  OAI2BB2XL U1676 ( .B0(n1457), .B1(n1514), .A0N(\gbuff[31][27] ), .A1N(n1515), 
        .Y(n1165) );
  OAI2BB2XL U1677 ( .B0(n1455), .B1(n1514), .A0N(\gbuff[31][28] ), .A1N(n1515), 
        .Y(n1166) );
  OAI2BB2XL U1678 ( .B0(n1453), .B1(n1514), .A0N(\gbuff[31][29] ), .A1N(n1515), 
        .Y(n1167) );
  OAI2BB2XL U1679 ( .B0(n1451), .B1(n1514), .A0N(\gbuff[31][30] ), .A1N(n1515), 
        .Y(n1168) );
  OAI2BB2XL U1680 ( .B0(n1449), .B1(n1514), .A0N(\gbuff[31][31] ), .A1N(n1513), 
        .Y(n1169) );
endmodule


module global_buffer_2 ( clk, rst, wr_en, index, data_in, data_out );
  input [7:0] index;
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, wr_en;
  wire   N10, N11, N12, N13, N14, \gbuff[1][31] , \gbuff[1][30] ,
         \gbuff[1][29] , \gbuff[1][28] , \gbuff[1][27] , \gbuff[1][26] ,
         \gbuff[1][25] , \gbuff[1][24] , \gbuff[1][23] , \gbuff[1][22] ,
         \gbuff[1][21] , \gbuff[1][20] , \gbuff[1][19] , \gbuff[1][18] ,
         \gbuff[1][17] , \gbuff[1][16] , \gbuff[1][15] , \gbuff[1][14] ,
         \gbuff[1][13] , \gbuff[1][12] , \gbuff[1][11] , \gbuff[1][10] ,
         \gbuff[1][9] , \gbuff[1][8] , \gbuff[1][7] , \gbuff[1][6] ,
         \gbuff[1][5] , \gbuff[1][4] , \gbuff[1][3] , \gbuff[1][2] ,
         \gbuff[1][1] , \gbuff[1][0] , \gbuff[0][31] , \gbuff[0][30] ,
         \gbuff[0][29] , \gbuff[0][28] , \gbuff[0][27] , \gbuff[0][26] ,
         \gbuff[0][25] , \gbuff[0][24] , \gbuff[0][23] , \gbuff[0][22] ,
         \gbuff[0][21] , \gbuff[0][20] , \gbuff[0][19] , \gbuff[0][18] ,
         \gbuff[0][17] , \gbuff[0][16] , \gbuff[0][15] , \gbuff[0][14] ,
         \gbuff[0][13] , \gbuff[0][12] , \gbuff[0][11] , \gbuff[0][10] ,
         \gbuff[0][9] , \gbuff[0][8] , \gbuff[0][7] , \gbuff[0][6] ,
         \gbuff[0][5] , \gbuff[0][4] , \gbuff[0][3] , \gbuff[0][2] ,
         \gbuff[0][1] , \gbuff[0][0] , \gbuff[3][31] , \gbuff[3][30] ,
         \gbuff[3][29] , \gbuff[3][28] , \gbuff[3][27] , \gbuff[3][26] ,
         \gbuff[3][25] , \gbuff[3][24] , \gbuff[3][23] , \gbuff[3][22] ,
         \gbuff[3][21] , \gbuff[3][20] , \gbuff[3][19] , \gbuff[3][18] ,
         \gbuff[3][17] , \gbuff[3][16] , \gbuff[3][15] , \gbuff[3][14] ,
         \gbuff[3][13] , \gbuff[3][12] , \gbuff[3][11] , \gbuff[3][10] ,
         \gbuff[3][9] , \gbuff[3][8] , \gbuff[3][7] , \gbuff[3][6] ,
         \gbuff[3][5] , \gbuff[3][4] , \gbuff[3][3] , \gbuff[3][2] ,
         \gbuff[3][1] , \gbuff[3][0] , \gbuff[2][31] , \gbuff[2][30] ,
         \gbuff[2][29] , \gbuff[2][28] , \gbuff[2][27] , \gbuff[2][26] ,
         \gbuff[2][25] , \gbuff[2][24] , \gbuff[2][23] , \gbuff[2][22] ,
         \gbuff[2][21] , \gbuff[2][20] , \gbuff[2][19] , \gbuff[2][18] ,
         \gbuff[2][17] , \gbuff[2][16] , \gbuff[2][15] , \gbuff[2][14] ,
         \gbuff[2][13] , \gbuff[2][12] , \gbuff[2][11] , \gbuff[2][10] ,
         \gbuff[2][9] , \gbuff[2][8] , \gbuff[2][7] , \gbuff[2][6] ,
         \gbuff[2][5] , \gbuff[2][4] , \gbuff[2][3] , \gbuff[2][2] ,
         \gbuff[2][1] , \gbuff[2][0] , \gbuff[5][31] , \gbuff[5][30] ,
         \gbuff[5][29] , \gbuff[5][28] , \gbuff[5][27] , \gbuff[5][26] ,
         \gbuff[5][25] , \gbuff[5][24] , \gbuff[5][23] , \gbuff[5][22] ,
         \gbuff[5][21] , \gbuff[5][20] , \gbuff[5][19] , \gbuff[5][18] ,
         \gbuff[5][17] , \gbuff[5][16] , \gbuff[5][15] , \gbuff[5][14] ,
         \gbuff[5][13] , \gbuff[5][12] , \gbuff[5][11] , \gbuff[5][10] ,
         \gbuff[5][9] , \gbuff[5][8] , \gbuff[5][7] , \gbuff[5][6] ,
         \gbuff[5][5] , \gbuff[5][4] , \gbuff[5][3] , \gbuff[5][2] ,
         \gbuff[5][1] , \gbuff[5][0] , \gbuff[4][31] , \gbuff[4][30] ,
         \gbuff[4][29] , \gbuff[4][28] , \gbuff[4][27] , \gbuff[4][26] ,
         \gbuff[4][25] , \gbuff[4][24] , \gbuff[4][23] , \gbuff[4][22] ,
         \gbuff[4][21] , \gbuff[4][20] , \gbuff[4][19] , \gbuff[4][18] ,
         \gbuff[4][17] , \gbuff[4][16] , \gbuff[4][15] , \gbuff[4][14] ,
         \gbuff[4][13] , \gbuff[4][12] , \gbuff[4][11] , \gbuff[4][10] ,
         \gbuff[4][9] , \gbuff[4][8] , \gbuff[4][7] , \gbuff[4][6] ,
         \gbuff[4][5] , \gbuff[4][4] , \gbuff[4][3] , \gbuff[4][2] ,
         \gbuff[4][1] , \gbuff[4][0] , \gbuff[7][31] , \gbuff[7][30] ,
         \gbuff[7][29] , \gbuff[7][28] , \gbuff[7][27] , \gbuff[7][26] ,
         \gbuff[7][25] , \gbuff[7][24] , \gbuff[7][23] , \gbuff[7][22] ,
         \gbuff[7][21] , \gbuff[7][20] , \gbuff[7][19] , \gbuff[7][18] ,
         \gbuff[7][17] , \gbuff[7][16] , \gbuff[7][15] , \gbuff[7][14] ,
         \gbuff[7][13] , \gbuff[7][12] , \gbuff[7][11] , \gbuff[7][10] ,
         \gbuff[7][9] , \gbuff[7][8] , \gbuff[7][7] , \gbuff[7][6] ,
         \gbuff[7][5] , \gbuff[7][4] , \gbuff[7][3] , \gbuff[7][2] ,
         \gbuff[7][1] , \gbuff[7][0] , \gbuff[6][31] , \gbuff[6][30] ,
         \gbuff[6][29] , \gbuff[6][28] , \gbuff[6][27] , \gbuff[6][26] ,
         \gbuff[6][25] , \gbuff[6][24] , \gbuff[6][23] , \gbuff[6][22] ,
         \gbuff[6][21] , \gbuff[6][20] , \gbuff[6][19] , \gbuff[6][18] ,
         \gbuff[6][17] , \gbuff[6][16] , \gbuff[6][15] , \gbuff[6][14] ,
         \gbuff[6][13] , \gbuff[6][12] , \gbuff[6][11] , \gbuff[6][10] ,
         \gbuff[6][9] , \gbuff[6][8] , \gbuff[6][7] , \gbuff[6][6] ,
         \gbuff[6][5] , \gbuff[6][4] , \gbuff[6][3] , \gbuff[6][2] ,
         \gbuff[6][1] , \gbuff[6][0] , \gbuff[9][31] , \gbuff[9][30] ,
         \gbuff[9][29] , \gbuff[9][28] , \gbuff[9][27] , \gbuff[9][26] ,
         \gbuff[9][25] , \gbuff[9][24] , \gbuff[9][23] , \gbuff[9][22] ,
         \gbuff[9][21] , \gbuff[9][20] , \gbuff[9][19] , \gbuff[9][18] ,
         \gbuff[9][17] , \gbuff[9][16] , \gbuff[9][15] , \gbuff[9][14] ,
         \gbuff[9][13] , \gbuff[9][12] , \gbuff[9][11] , \gbuff[9][10] ,
         \gbuff[9][9] , \gbuff[9][8] , \gbuff[9][7] , \gbuff[9][6] ,
         \gbuff[9][5] , \gbuff[9][4] , \gbuff[9][3] , \gbuff[9][2] ,
         \gbuff[9][1] , \gbuff[9][0] , \gbuff[8][31] , \gbuff[8][30] ,
         \gbuff[8][29] , \gbuff[8][28] , \gbuff[8][27] , \gbuff[8][26] ,
         \gbuff[8][25] , \gbuff[8][24] , \gbuff[8][23] , \gbuff[8][22] ,
         \gbuff[8][21] , \gbuff[8][20] , \gbuff[8][19] , \gbuff[8][18] ,
         \gbuff[8][17] , \gbuff[8][16] , \gbuff[8][15] , \gbuff[8][14] ,
         \gbuff[8][13] , \gbuff[8][12] , \gbuff[8][11] , \gbuff[8][10] ,
         \gbuff[8][9] , \gbuff[8][8] , \gbuff[8][7] , \gbuff[8][6] ,
         \gbuff[8][5] , \gbuff[8][4] , \gbuff[8][3] , \gbuff[8][2] ,
         \gbuff[8][1] , \gbuff[8][0] , \gbuff[11][31] , \gbuff[11][30] ,
         \gbuff[11][29] , \gbuff[11][28] , \gbuff[11][27] , \gbuff[11][26] ,
         \gbuff[11][25] , \gbuff[11][24] , \gbuff[11][23] , \gbuff[11][22] ,
         \gbuff[11][21] , \gbuff[11][20] , \gbuff[11][19] , \gbuff[11][18] ,
         \gbuff[11][17] , \gbuff[11][16] , \gbuff[11][15] , \gbuff[11][14] ,
         \gbuff[11][13] , \gbuff[11][12] , \gbuff[11][11] , \gbuff[11][10] ,
         \gbuff[11][9] , \gbuff[11][8] , \gbuff[11][7] , \gbuff[11][6] ,
         \gbuff[11][5] , \gbuff[11][4] , \gbuff[11][3] , \gbuff[11][2] ,
         \gbuff[11][1] , \gbuff[11][0] , \gbuff[10][31] , \gbuff[10][30] ,
         \gbuff[10][29] , \gbuff[10][28] , \gbuff[10][27] , \gbuff[10][26] ,
         \gbuff[10][25] , \gbuff[10][24] , \gbuff[10][23] , \gbuff[10][22] ,
         \gbuff[10][21] , \gbuff[10][20] , \gbuff[10][19] , \gbuff[10][18] ,
         \gbuff[10][17] , \gbuff[10][16] , \gbuff[10][15] , \gbuff[10][14] ,
         \gbuff[10][13] , \gbuff[10][12] , \gbuff[10][11] , \gbuff[10][10] ,
         \gbuff[10][9] , \gbuff[10][8] , \gbuff[10][7] , \gbuff[10][6] ,
         \gbuff[10][5] , \gbuff[10][4] , \gbuff[10][3] , \gbuff[10][2] ,
         \gbuff[10][1] , \gbuff[10][0] , \gbuff[13][31] , \gbuff[13][30] ,
         \gbuff[13][29] , \gbuff[13][28] , \gbuff[13][27] , \gbuff[13][26] ,
         \gbuff[13][25] , \gbuff[13][24] , \gbuff[13][23] , \gbuff[13][22] ,
         \gbuff[13][21] , \gbuff[13][20] , \gbuff[13][19] , \gbuff[13][18] ,
         \gbuff[13][17] , \gbuff[13][16] , \gbuff[13][15] , \gbuff[13][14] ,
         \gbuff[13][13] , \gbuff[13][12] , \gbuff[13][11] , \gbuff[13][10] ,
         \gbuff[13][9] , \gbuff[13][8] , \gbuff[13][7] , \gbuff[13][6] ,
         \gbuff[13][5] , \gbuff[13][4] , \gbuff[13][3] , \gbuff[13][2] ,
         \gbuff[13][1] , \gbuff[13][0] , \gbuff[12][31] , \gbuff[12][30] ,
         \gbuff[12][29] , \gbuff[12][28] , \gbuff[12][27] , \gbuff[12][26] ,
         \gbuff[12][25] , \gbuff[12][24] , \gbuff[12][23] , \gbuff[12][22] ,
         \gbuff[12][21] , \gbuff[12][20] , \gbuff[12][19] , \gbuff[12][18] ,
         \gbuff[12][17] , \gbuff[12][16] , \gbuff[12][15] , \gbuff[12][14] ,
         \gbuff[12][13] , \gbuff[12][12] , \gbuff[12][11] , \gbuff[12][10] ,
         \gbuff[12][9] , \gbuff[12][8] , \gbuff[12][7] , \gbuff[12][6] ,
         \gbuff[12][5] , \gbuff[12][4] , \gbuff[12][3] , \gbuff[12][2] ,
         \gbuff[12][1] , \gbuff[12][0] , \gbuff[15][31] , \gbuff[15][30] ,
         \gbuff[15][29] , \gbuff[15][28] , \gbuff[15][27] , \gbuff[15][26] ,
         \gbuff[15][25] , \gbuff[15][24] , \gbuff[15][23] , \gbuff[15][22] ,
         \gbuff[15][21] , \gbuff[15][20] , \gbuff[15][19] , \gbuff[15][18] ,
         \gbuff[15][17] , \gbuff[15][16] , \gbuff[15][15] , \gbuff[15][14] ,
         \gbuff[15][13] , \gbuff[15][12] , \gbuff[15][11] , \gbuff[15][10] ,
         \gbuff[15][9] , \gbuff[15][8] , \gbuff[15][7] , \gbuff[15][6] ,
         \gbuff[15][5] , \gbuff[15][4] , \gbuff[15][3] , \gbuff[15][2] ,
         \gbuff[15][1] , \gbuff[15][0] , \gbuff[14][31] , \gbuff[14][30] ,
         \gbuff[14][29] , \gbuff[14][28] , \gbuff[14][27] , \gbuff[14][26] ,
         \gbuff[14][25] , \gbuff[14][24] , \gbuff[14][23] , \gbuff[14][22] ,
         \gbuff[14][21] , \gbuff[14][20] , \gbuff[14][19] , \gbuff[14][18] ,
         \gbuff[14][17] , \gbuff[14][16] , \gbuff[14][15] , \gbuff[14][14] ,
         \gbuff[14][13] , \gbuff[14][12] , \gbuff[14][11] , \gbuff[14][10] ,
         \gbuff[14][9] , \gbuff[14][8] , \gbuff[14][7] , \gbuff[14][6] ,
         \gbuff[14][5] , \gbuff[14][4] , \gbuff[14][3] , \gbuff[14][2] ,
         \gbuff[14][1] , \gbuff[14][0] , \gbuff[17][31] , \gbuff[17][30] ,
         \gbuff[17][29] , \gbuff[17][28] , \gbuff[17][27] , \gbuff[17][26] ,
         \gbuff[17][25] , \gbuff[17][24] , \gbuff[17][23] , \gbuff[17][22] ,
         \gbuff[17][21] , \gbuff[17][20] , \gbuff[17][19] , \gbuff[17][18] ,
         \gbuff[17][17] , \gbuff[17][16] , \gbuff[17][15] , \gbuff[17][14] ,
         \gbuff[17][13] , \gbuff[17][12] , \gbuff[17][11] , \gbuff[17][10] ,
         \gbuff[17][9] , \gbuff[17][8] , \gbuff[17][7] , \gbuff[17][6] ,
         \gbuff[17][5] , \gbuff[17][4] , \gbuff[17][3] , \gbuff[17][2] ,
         \gbuff[17][1] , \gbuff[17][0] , \gbuff[16][31] , \gbuff[16][30] ,
         \gbuff[16][29] , \gbuff[16][28] , \gbuff[16][27] , \gbuff[16][26] ,
         \gbuff[16][25] , \gbuff[16][24] , \gbuff[16][23] , \gbuff[16][22] ,
         \gbuff[16][21] , \gbuff[16][20] , \gbuff[16][19] , \gbuff[16][18] ,
         \gbuff[16][17] , \gbuff[16][16] , \gbuff[16][15] , \gbuff[16][14] ,
         \gbuff[16][13] , \gbuff[16][12] , \gbuff[16][11] , \gbuff[16][10] ,
         \gbuff[16][9] , \gbuff[16][8] , \gbuff[16][7] , \gbuff[16][6] ,
         \gbuff[16][5] , \gbuff[16][4] , \gbuff[16][3] , \gbuff[16][2] ,
         \gbuff[16][1] , \gbuff[16][0] , \gbuff[19][31] , \gbuff[19][30] ,
         \gbuff[19][29] , \gbuff[19][28] , \gbuff[19][27] , \gbuff[19][26] ,
         \gbuff[19][25] , \gbuff[19][24] , \gbuff[19][23] , \gbuff[19][22] ,
         \gbuff[19][21] , \gbuff[19][20] , \gbuff[19][19] , \gbuff[19][18] ,
         \gbuff[19][17] , \gbuff[19][16] , \gbuff[19][15] , \gbuff[19][14] ,
         \gbuff[19][13] , \gbuff[19][12] , \gbuff[19][11] , \gbuff[19][10] ,
         \gbuff[19][9] , \gbuff[19][8] , \gbuff[19][7] , \gbuff[19][6] ,
         \gbuff[19][5] , \gbuff[19][4] , \gbuff[19][3] , \gbuff[19][2] ,
         \gbuff[19][1] , \gbuff[19][0] , \gbuff[18][31] , \gbuff[18][30] ,
         \gbuff[18][29] , \gbuff[18][28] , \gbuff[18][27] , \gbuff[18][26] ,
         \gbuff[18][25] , \gbuff[18][24] , \gbuff[18][23] , \gbuff[18][22] ,
         \gbuff[18][21] , \gbuff[18][20] , \gbuff[18][19] , \gbuff[18][18] ,
         \gbuff[18][17] , \gbuff[18][16] , \gbuff[18][15] , \gbuff[18][14] ,
         \gbuff[18][13] , \gbuff[18][12] , \gbuff[18][11] , \gbuff[18][10] ,
         \gbuff[18][9] , \gbuff[18][8] , \gbuff[18][7] , \gbuff[18][6] ,
         \gbuff[18][5] , \gbuff[18][4] , \gbuff[18][3] , \gbuff[18][2] ,
         \gbuff[18][1] , \gbuff[18][0] , \gbuff[21][31] , \gbuff[21][30] ,
         \gbuff[21][29] , \gbuff[21][28] , \gbuff[21][27] , \gbuff[21][26] ,
         \gbuff[21][25] , \gbuff[21][24] , \gbuff[21][23] , \gbuff[21][22] ,
         \gbuff[21][21] , \gbuff[21][20] , \gbuff[21][19] , \gbuff[21][18] ,
         \gbuff[21][17] , \gbuff[21][16] , \gbuff[21][15] , \gbuff[21][14] ,
         \gbuff[21][13] , \gbuff[21][12] , \gbuff[21][11] , \gbuff[21][10] ,
         \gbuff[21][9] , \gbuff[21][8] , \gbuff[21][7] , \gbuff[21][6] ,
         \gbuff[21][5] , \gbuff[21][4] , \gbuff[21][3] , \gbuff[21][2] ,
         \gbuff[21][1] , \gbuff[21][0] , \gbuff[20][31] , \gbuff[20][30] ,
         \gbuff[20][29] , \gbuff[20][28] , \gbuff[20][27] , \gbuff[20][26] ,
         \gbuff[20][25] , \gbuff[20][24] , \gbuff[20][23] , \gbuff[20][22] ,
         \gbuff[20][21] , \gbuff[20][20] , \gbuff[20][19] , \gbuff[20][18] ,
         \gbuff[20][17] , \gbuff[20][16] , \gbuff[20][15] , \gbuff[20][14] ,
         \gbuff[20][13] , \gbuff[20][12] , \gbuff[20][11] , \gbuff[20][10] ,
         \gbuff[20][9] , \gbuff[20][8] , \gbuff[20][7] , \gbuff[20][6] ,
         \gbuff[20][5] , \gbuff[20][4] , \gbuff[20][3] , \gbuff[20][2] ,
         \gbuff[20][1] , \gbuff[20][0] , \gbuff[23][31] , \gbuff[23][30] ,
         \gbuff[23][29] , \gbuff[23][28] , \gbuff[23][27] , \gbuff[23][26] ,
         \gbuff[23][25] , \gbuff[23][24] , \gbuff[23][23] , \gbuff[23][22] ,
         \gbuff[23][21] , \gbuff[23][20] , \gbuff[23][19] , \gbuff[23][18] ,
         \gbuff[23][17] , \gbuff[23][16] , \gbuff[23][15] , \gbuff[23][14] ,
         \gbuff[23][13] , \gbuff[23][12] , \gbuff[23][11] , \gbuff[23][10] ,
         \gbuff[23][9] , \gbuff[23][8] , \gbuff[23][7] , \gbuff[23][6] ,
         \gbuff[23][5] , \gbuff[23][4] , \gbuff[23][3] , \gbuff[23][2] ,
         \gbuff[23][1] , \gbuff[23][0] , \gbuff[22][31] , \gbuff[22][30] ,
         \gbuff[22][29] , \gbuff[22][28] , \gbuff[22][27] , \gbuff[22][26] ,
         \gbuff[22][25] , \gbuff[22][24] , \gbuff[22][23] , \gbuff[22][22] ,
         \gbuff[22][21] , \gbuff[22][20] , \gbuff[22][19] , \gbuff[22][18] ,
         \gbuff[22][17] , \gbuff[22][16] , \gbuff[22][15] , \gbuff[22][14] ,
         \gbuff[22][13] , \gbuff[22][12] , \gbuff[22][11] , \gbuff[22][10] ,
         \gbuff[22][9] , \gbuff[22][8] , \gbuff[22][7] , \gbuff[22][6] ,
         \gbuff[22][5] , \gbuff[22][4] , \gbuff[22][3] , \gbuff[22][2] ,
         \gbuff[22][1] , \gbuff[22][0] , \gbuff[25][31] , \gbuff[25][30] ,
         \gbuff[25][29] , \gbuff[25][28] , \gbuff[25][27] , \gbuff[25][26] ,
         \gbuff[25][25] , \gbuff[25][24] , \gbuff[25][23] , \gbuff[25][22] ,
         \gbuff[25][21] , \gbuff[25][20] , \gbuff[25][19] , \gbuff[25][18] ,
         \gbuff[25][17] , \gbuff[25][16] , \gbuff[25][15] , \gbuff[25][14] ,
         \gbuff[25][13] , \gbuff[25][12] , \gbuff[25][11] , \gbuff[25][10] ,
         \gbuff[25][9] , \gbuff[25][8] , \gbuff[25][7] , \gbuff[25][6] ,
         \gbuff[25][5] , \gbuff[25][4] , \gbuff[25][3] , \gbuff[25][2] ,
         \gbuff[25][1] , \gbuff[25][0] , \gbuff[24][31] , \gbuff[24][30] ,
         \gbuff[24][29] , \gbuff[24][28] , \gbuff[24][27] , \gbuff[24][26] ,
         \gbuff[24][25] , \gbuff[24][24] , \gbuff[24][23] , \gbuff[24][22] ,
         \gbuff[24][21] , \gbuff[24][20] , \gbuff[24][19] , \gbuff[24][18] ,
         \gbuff[24][17] , \gbuff[24][16] , \gbuff[24][15] , \gbuff[24][14] ,
         \gbuff[24][13] , \gbuff[24][12] , \gbuff[24][11] , \gbuff[24][10] ,
         \gbuff[24][9] , \gbuff[24][8] , \gbuff[24][7] , \gbuff[24][6] ,
         \gbuff[24][5] , \gbuff[24][4] , \gbuff[24][3] , \gbuff[24][2] ,
         \gbuff[24][1] , \gbuff[24][0] , \gbuff[27][31] , \gbuff[27][30] ,
         \gbuff[27][29] , \gbuff[27][28] , \gbuff[27][27] , \gbuff[27][26] ,
         \gbuff[27][25] , \gbuff[27][24] , \gbuff[27][23] , \gbuff[27][22] ,
         \gbuff[27][21] , \gbuff[27][20] , \gbuff[27][19] , \gbuff[27][18] ,
         \gbuff[27][17] , \gbuff[27][16] , \gbuff[27][15] , \gbuff[27][14] ,
         \gbuff[27][13] , \gbuff[27][12] , \gbuff[27][11] , \gbuff[27][10] ,
         \gbuff[27][9] , \gbuff[27][8] , \gbuff[27][7] , \gbuff[27][6] ,
         \gbuff[27][5] , \gbuff[27][4] , \gbuff[27][3] , \gbuff[27][2] ,
         \gbuff[27][1] , \gbuff[27][0] , \gbuff[26][31] , \gbuff[26][30] ,
         \gbuff[26][29] , \gbuff[26][28] , \gbuff[26][27] , \gbuff[26][26] ,
         \gbuff[26][25] , \gbuff[26][24] , \gbuff[26][23] , \gbuff[26][22] ,
         \gbuff[26][21] , \gbuff[26][20] , \gbuff[26][19] , \gbuff[26][18] ,
         \gbuff[26][17] , \gbuff[26][16] , \gbuff[26][15] , \gbuff[26][14] ,
         \gbuff[26][13] , \gbuff[26][12] , \gbuff[26][11] , \gbuff[26][10] ,
         \gbuff[26][9] , \gbuff[26][8] , \gbuff[26][7] , \gbuff[26][6] ,
         \gbuff[26][5] , \gbuff[26][4] , \gbuff[26][3] , \gbuff[26][2] ,
         \gbuff[26][1] , \gbuff[26][0] , \gbuff[29][31] , \gbuff[29][30] ,
         \gbuff[29][29] , \gbuff[29][28] , \gbuff[29][27] , \gbuff[29][26] ,
         \gbuff[29][25] , \gbuff[29][24] , \gbuff[29][23] , \gbuff[29][22] ,
         \gbuff[29][21] , \gbuff[29][20] , \gbuff[29][19] , \gbuff[29][18] ,
         \gbuff[29][17] , \gbuff[29][16] , \gbuff[29][15] , \gbuff[29][14] ,
         \gbuff[29][13] , \gbuff[29][12] , \gbuff[29][11] , \gbuff[29][10] ,
         \gbuff[29][9] , \gbuff[29][8] , \gbuff[29][7] , \gbuff[29][6] ,
         \gbuff[29][5] , \gbuff[29][4] , \gbuff[29][3] , \gbuff[29][2] ,
         \gbuff[29][1] , \gbuff[29][0] , \gbuff[28][31] , \gbuff[28][30] ,
         \gbuff[28][29] , \gbuff[28][28] , \gbuff[28][27] , \gbuff[28][26] ,
         \gbuff[28][25] , \gbuff[28][24] , \gbuff[28][23] , \gbuff[28][22] ,
         \gbuff[28][21] , \gbuff[28][20] , \gbuff[28][19] , \gbuff[28][18] ,
         \gbuff[28][17] , \gbuff[28][16] , \gbuff[28][15] , \gbuff[28][14] ,
         \gbuff[28][13] , \gbuff[28][12] , \gbuff[28][11] , \gbuff[28][10] ,
         \gbuff[28][9] , \gbuff[28][8] , \gbuff[28][7] , \gbuff[28][6] ,
         \gbuff[28][5] , \gbuff[28][4] , \gbuff[28][3] , \gbuff[28][2] ,
         \gbuff[28][1] , \gbuff[28][0] , \gbuff[31][31] , \gbuff[31][30] ,
         \gbuff[31][29] , \gbuff[31][28] , \gbuff[31][27] , \gbuff[31][26] ,
         \gbuff[31][25] , \gbuff[31][24] , \gbuff[31][23] , \gbuff[31][22] ,
         \gbuff[31][21] , \gbuff[31][20] , \gbuff[31][19] , \gbuff[31][18] ,
         \gbuff[31][17] , \gbuff[31][16] , \gbuff[31][15] , \gbuff[31][14] ,
         \gbuff[31][13] , \gbuff[31][12] , \gbuff[31][11] , \gbuff[31][10] ,
         \gbuff[31][9] , \gbuff[31][8] , \gbuff[31][7] , \gbuff[31][6] ,
         \gbuff[31][5] , \gbuff[31][4] , \gbuff[31][3] , \gbuff[31][2] ,
         \gbuff[31][1] , \gbuff[31][0] , \gbuff[30][31] , \gbuff[30][30] ,
         \gbuff[30][29] , \gbuff[30][28] , \gbuff[30][27] , \gbuff[30][26] ,
         \gbuff[30][25] , \gbuff[30][24] , \gbuff[30][23] , \gbuff[30][22] ,
         \gbuff[30][21] , \gbuff[30][20] , \gbuff[30][19] , \gbuff[30][18] ,
         \gbuff[30][17] , \gbuff[30][16] , \gbuff[30][15] , \gbuff[30][14] ,
         \gbuff[30][13] , \gbuff[30][12] , \gbuff[30][11] , \gbuff[30][10] ,
         \gbuff[30][9] , \gbuff[30][8] , \gbuff[30][7] , \gbuff[30][6] ,
         \gbuff[30][5] , \gbuff[30][4] , \gbuff[30][3] , \gbuff[30][2] ,
         \gbuff[30][1] , \gbuff[30][0] , N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N81, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n104,
         n106, n108, n110, n112, n114, n116, n119, n121, n122, n123, n124,
         n125, n126, n127, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847;
  assign N10 = index[0];
  assign N11 = index[1];
  assign N12 = index[2];
  assign N13 = index[3];
  assign N14 = index[4];

  DFFRX1 \gbuff_reg[29][31]  ( .D(n1859), .CK(clk), .RN(n1601), .Q(
        \gbuff[29][31] ) );
  DFFRX1 \gbuff_reg[29][30]  ( .D(n1860), .CK(clk), .RN(n1601), .Q(
        \gbuff[29][30] ) );
  DFFRX1 \gbuff_reg[29][29]  ( .D(n1861), .CK(clk), .RN(n1601), .Q(
        \gbuff[29][29] ) );
  DFFRX1 \gbuff_reg[29][28]  ( .D(n1862), .CK(clk), .RN(n1601), .Q(
        \gbuff[29][28] ) );
  DFFRX1 \gbuff_reg[29][27]  ( .D(n1863), .CK(clk), .RN(n1601), .Q(
        \gbuff[29][27] ) );
  DFFRX1 \gbuff_reg[29][26]  ( .D(n1864), .CK(clk), .RN(n1601), .Q(
        \gbuff[29][26] ) );
  DFFRX1 \gbuff_reg[29][25]  ( .D(n1865), .CK(clk), .RN(n1601), .Q(
        \gbuff[29][25] ) );
  DFFRX1 \gbuff_reg[29][24]  ( .D(n1866), .CK(clk), .RN(n1601), .Q(
        \gbuff[29][24] ) );
  DFFRX1 \gbuff_reg[29][23]  ( .D(n1867), .CK(clk), .RN(n1601), .Q(
        \gbuff[29][23] ) );
  DFFRX1 \gbuff_reg[29][22]  ( .D(n1868), .CK(clk), .RN(n1601), .Q(
        \gbuff[29][22] ) );
  DFFRX1 \gbuff_reg[29][21]  ( .D(n1869), .CK(clk), .RN(n1601), .Q(
        \gbuff[29][21] ) );
  DFFRX1 \gbuff_reg[29][20]  ( .D(n1870), .CK(clk), .RN(n1601), .Q(
        \gbuff[29][20] ) );
  DFFRX1 \gbuff_reg[29][19]  ( .D(n1871), .CK(clk), .RN(n1600), .Q(
        \gbuff[29][19] ) );
  DFFRX1 \gbuff_reg[29][18]  ( .D(n1872), .CK(clk), .RN(n1600), .Q(
        \gbuff[29][18] ) );
  DFFRX1 \gbuff_reg[29][17]  ( .D(n1873), .CK(clk), .RN(n1600), .Q(
        \gbuff[29][17] ) );
  DFFRX1 \gbuff_reg[29][16]  ( .D(n1874), .CK(clk), .RN(n1600), .Q(
        \gbuff[29][16] ) );
  DFFRX1 \gbuff_reg[29][15]  ( .D(n1875), .CK(clk), .RN(n1600), .Q(
        \gbuff[29][15] ) );
  DFFRX1 \gbuff_reg[29][14]  ( .D(n1876), .CK(clk), .RN(n1600), .Q(
        \gbuff[29][14] ) );
  DFFRX1 \gbuff_reg[29][13]  ( .D(n1877), .CK(clk), .RN(n1600), .Q(
        \gbuff[29][13] ) );
  DFFRX1 \gbuff_reg[29][12]  ( .D(n1878), .CK(clk), .RN(n1600), .Q(
        \gbuff[29][12] ) );
  DFFRX1 \gbuff_reg[29][11]  ( .D(n1879), .CK(clk), .RN(n1600), .Q(
        \gbuff[29][11] ) );
  DFFRX1 \gbuff_reg[29][10]  ( .D(n1880), .CK(clk), .RN(n1600), .Q(
        \gbuff[29][10] ) );
  DFFRX1 \gbuff_reg[29][9]  ( .D(n1881), .CK(clk), .RN(n1600), .Q(
        \gbuff[29][9] ) );
  DFFRX1 \gbuff_reg[29][8]  ( .D(n1882), .CK(clk), .RN(n1600), .Q(
        \gbuff[29][8] ) );
  DFFRX1 \gbuff_reg[29][7]  ( .D(n1883), .CK(clk), .RN(n1599), .Q(
        \gbuff[29][7] ) );
  DFFRX1 \gbuff_reg[29][6]  ( .D(n1884), .CK(clk), .RN(n1599), .Q(
        \gbuff[29][6] ) );
  DFFRX1 \gbuff_reg[29][5]  ( .D(n1885), .CK(clk), .RN(n1599), .Q(
        \gbuff[29][5] ) );
  DFFRX1 \gbuff_reg[29][4]  ( .D(n1886), .CK(clk), .RN(n1599), .Q(
        \gbuff[29][4] ) );
  DFFRX1 \gbuff_reg[29][3]  ( .D(n1887), .CK(clk), .RN(n1599), .Q(
        \gbuff[29][3] ) );
  DFFRX1 \gbuff_reg[29][2]  ( .D(n1888), .CK(clk), .RN(n1599), .Q(
        \gbuff[29][2] ) );
  DFFRX1 \gbuff_reg[29][1]  ( .D(n1889), .CK(clk), .RN(n1599), .Q(
        \gbuff[29][1] ) );
  DFFRX1 \gbuff_reg[29][0]  ( .D(n1890), .CK(clk), .RN(n1599), .Q(
        \gbuff[29][0] ) );
  DFFRX1 \gbuff_reg[25][31]  ( .D(n1987), .CK(clk), .RN(n1591), .Q(
        \gbuff[25][31] ) );
  DFFRX1 \gbuff_reg[25][30]  ( .D(n1988), .CK(clk), .RN(n1591), .Q(
        \gbuff[25][30] ) );
  DFFRX1 \gbuff_reg[25][29]  ( .D(n1989), .CK(clk), .RN(n1591), .Q(
        \gbuff[25][29] ) );
  DFFRX1 \gbuff_reg[25][28]  ( .D(n1990), .CK(clk), .RN(n1591), .Q(
        \gbuff[25][28] ) );
  DFFRX1 \gbuff_reg[25][27]  ( .D(n1991), .CK(clk), .RN(n1590), .Q(
        \gbuff[25][27] ) );
  DFFRX1 \gbuff_reg[25][26]  ( .D(n1992), .CK(clk), .RN(n1590), .Q(
        \gbuff[25][26] ) );
  DFFRX1 \gbuff_reg[25][25]  ( .D(n1993), .CK(clk), .RN(n1590), .Q(
        \gbuff[25][25] ) );
  DFFRX1 \gbuff_reg[25][24]  ( .D(n1994), .CK(clk), .RN(n1590), .Q(
        \gbuff[25][24] ) );
  DFFRX1 \gbuff_reg[25][23]  ( .D(n1995), .CK(clk), .RN(n1590), .Q(
        \gbuff[25][23] ) );
  DFFRX1 \gbuff_reg[25][22]  ( .D(n1996), .CK(clk), .RN(n1590), .Q(
        \gbuff[25][22] ) );
  DFFRX1 \gbuff_reg[25][21]  ( .D(n1997), .CK(clk), .RN(n1590), .Q(
        \gbuff[25][21] ) );
  DFFRX1 \gbuff_reg[25][20]  ( .D(n1998), .CK(clk), .RN(n1590), .Q(
        \gbuff[25][20] ) );
  DFFRX1 \gbuff_reg[25][19]  ( .D(n1999), .CK(clk), .RN(n1590), .Q(
        \gbuff[25][19] ) );
  DFFRX1 \gbuff_reg[25][18]  ( .D(n2000), .CK(clk), .RN(n1590), .Q(
        \gbuff[25][18] ) );
  DFFRX1 \gbuff_reg[25][17]  ( .D(n2001), .CK(clk), .RN(n1590), .Q(
        \gbuff[25][17] ) );
  DFFRX1 \gbuff_reg[25][16]  ( .D(n2002), .CK(clk), .RN(n1590), .Q(
        \gbuff[25][16] ) );
  DFFRX1 \gbuff_reg[25][15]  ( .D(n2003), .CK(clk), .RN(n1589), .Q(
        \gbuff[25][15] ) );
  DFFRX1 \gbuff_reg[25][14]  ( .D(n2004), .CK(clk), .RN(n1589), .Q(
        \gbuff[25][14] ) );
  DFFRX1 \gbuff_reg[25][13]  ( .D(n2005), .CK(clk), .RN(n1589), .Q(
        \gbuff[25][13] ) );
  DFFRX1 \gbuff_reg[25][12]  ( .D(n2006), .CK(clk), .RN(n1589), .Q(
        \gbuff[25][12] ) );
  DFFRX1 \gbuff_reg[25][11]  ( .D(n2007), .CK(clk), .RN(n1589), .Q(
        \gbuff[25][11] ) );
  DFFRX1 \gbuff_reg[25][10]  ( .D(n2008), .CK(clk), .RN(n1589), .Q(
        \gbuff[25][10] ) );
  DFFRX1 \gbuff_reg[25][9]  ( .D(n2009), .CK(clk), .RN(n1589), .Q(
        \gbuff[25][9] ) );
  DFFRX1 \gbuff_reg[25][8]  ( .D(n2010), .CK(clk), .RN(n1589), .Q(
        \gbuff[25][8] ) );
  DFFRX1 \gbuff_reg[25][7]  ( .D(n2011), .CK(clk), .RN(n1589), .Q(
        \gbuff[25][7] ) );
  DFFRX1 \gbuff_reg[25][6]  ( .D(n2012), .CK(clk), .RN(n1589), .Q(
        \gbuff[25][6] ) );
  DFFRX1 \gbuff_reg[25][5]  ( .D(n2013), .CK(clk), .RN(n1589), .Q(
        \gbuff[25][5] ) );
  DFFRX1 \gbuff_reg[25][4]  ( .D(n2014), .CK(clk), .RN(n1589), .Q(
        \gbuff[25][4] ) );
  DFFRX1 \gbuff_reg[25][3]  ( .D(n2015), .CK(clk), .RN(n1588), .Q(
        \gbuff[25][3] ) );
  DFFRX1 \gbuff_reg[25][2]  ( .D(n2016), .CK(clk), .RN(n1588), .Q(
        \gbuff[25][2] ) );
  DFFRX1 \gbuff_reg[25][1]  ( .D(n2017), .CK(clk), .RN(n1588), .Q(
        \gbuff[25][1] ) );
  DFFRX1 \gbuff_reg[25][0]  ( .D(n2018), .CK(clk), .RN(n1588), .Q(
        \gbuff[25][0] ) );
  DFFRX1 \gbuff_reg[21][31]  ( .D(n2115), .CK(clk), .RN(n1580), .Q(
        \gbuff[21][31] ) );
  DFFRX1 \gbuff_reg[21][30]  ( .D(n2116), .CK(clk), .RN(n1580), .Q(
        \gbuff[21][30] ) );
  DFFRX1 \gbuff_reg[21][29]  ( .D(n2117), .CK(clk), .RN(n1580), .Q(
        \gbuff[21][29] ) );
  DFFRX1 \gbuff_reg[21][28]  ( .D(n2118), .CK(clk), .RN(n1580), .Q(
        \gbuff[21][28] ) );
  DFFRX1 \gbuff_reg[21][27]  ( .D(n2119), .CK(clk), .RN(n1580), .Q(
        \gbuff[21][27] ) );
  DFFRX1 \gbuff_reg[21][26]  ( .D(n2120), .CK(clk), .RN(n1580), .Q(
        \gbuff[21][26] ) );
  DFFRX1 \gbuff_reg[21][25]  ( .D(n2121), .CK(clk), .RN(n1580), .Q(
        \gbuff[21][25] ) );
  DFFRX1 \gbuff_reg[21][24]  ( .D(n2122), .CK(clk), .RN(n1580), .Q(
        \gbuff[21][24] ) );
  DFFRX1 \gbuff_reg[21][23]  ( .D(n2123), .CK(clk), .RN(n1579), .Q(
        \gbuff[21][23] ) );
  DFFRX1 \gbuff_reg[21][22]  ( .D(n2124), .CK(clk), .RN(n1579), .Q(
        \gbuff[21][22] ) );
  DFFRX1 \gbuff_reg[21][21]  ( .D(n2125), .CK(clk), .RN(n1579), .Q(
        \gbuff[21][21] ) );
  DFFRX1 \gbuff_reg[21][20]  ( .D(n2126), .CK(clk), .RN(n1579), .Q(
        \gbuff[21][20] ) );
  DFFRX1 \gbuff_reg[21][19]  ( .D(n2127), .CK(clk), .RN(n1579), .Q(
        \gbuff[21][19] ) );
  DFFRX1 \gbuff_reg[21][18]  ( .D(n2128), .CK(clk), .RN(n1579), .Q(
        \gbuff[21][18] ) );
  DFFRX1 \gbuff_reg[21][17]  ( .D(n2129), .CK(clk), .RN(n1579), .Q(
        \gbuff[21][17] ) );
  DFFRX1 \gbuff_reg[21][16]  ( .D(n2130), .CK(clk), .RN(n1579), .Q(
        \gbuff[21][16] ) );
  DFFRX1 \gbuff_reg[21][15]  ( .D(n2131), .CK(clk), .RN(n1579), .Q(
        \gbuff[21][15] ) );
  DFFRX1 \gbuff_reg[21][14]  ( .D(n2132), .CK(clk), .RN(n1579), .Q(
        \gbuff[21][14] ) );
  DFFRX1 \gbuff_reg[21][13]  ( .D(n2133), .CK(clk), .RN(n1579), .Q(
        \gbuff[21][13] ) );
  DFFRX1 \gbuff_reg[21][12]  ( .D(n2134), .CK(clk), .RN(n1579), .Q(
        \gbuff[21][12] ) );
  DFFRX1 \gbuff_reg[21][11]  ( .D(n2135), .CK(clk), .RN(n1578), .Q(
        \gbuff[21][11] ) );
  DFFRX1 \gbuff_reg[21][10]  ( .D(n2136), .CK(clk), .RN(n1578), .Q(
        \gbuff[21][10] ) );
  DFFRX1 \gbuff_reg[21][9]  ( .D(n2137), .CK(clk), .RN(n1578), .Q(
        \gbuff[21][9] ) );
  DFFRX1 \gbuff_reg[21][8]  ( .D(n2138), .CK(clk), .RN(n1578), .Q(
        \gbuff[21][8] ) );
  DFFRX1 \gbuff_reg[21][7]  ( .D(n2139), .CK(clk), .RN(n1578), .Q(
        \gbuff[21][7] ) );
  DFFRX1 \gbuff_reg[21][6]  ( .D(n2140), .CK(clk), .RN(n1578), .Q(
        \gbuff[21][6] ) );
  DFFRX1 \gbuff_reg[21][5]  ( .D(n2141), .CK(clk), .RN(n1578), .Q(
        \gbuff[21][5] ) );
  DFFRX1 \gbuff_reg[21][4]  ( .D(n2142), .CK(clk), .RN(n1578), .Q(
        \gbuff[21][4] ) );
  DFFRX1 \gbuff_reg[21][3]  ( .D(n2143), .CK(clk), .RN(n1578), .Q(
        \gbuff[21][3] ) );
  DFFRX1 \gbuff_reg[21][2]  ( .D(n2144), .CK(clk), .RN(n1578), .Q(
        \gbuff[21][2] ) );
  DFFRX1 \gbuff_reg[21][1]  ( .D(n2145), .CK(clk), .RN(n1578), .Q(
        \gbuff[21][1] ) );
  DFFRX1 \gbuff_reg[21][0]  ( .D(n2146), .CK(clk), .RN(n1578), .Q(
        \gbuff[21][0] ) );
  DFFRX1 \gbuff_reg[17][31]  ( .D(n2243), .CK(clk), .RN(n1569), .Q(
        \gbuff[17][31] ) );
  DFFRX1 \gbuff_reg[17][30]  ( .D(n2244), .CK(clk), .RN(n1569), .Q(
        \gbuff[17][30] ) );
  DFFRX1 \gbuff_reg[17][29]  ( .D(n2245), .CK(clk), .RN(n1569), .Q(
        \gbuff[17][29] ) );
  DFFRX1 \gbuff_reg[17][28]  ( .D(n2246), .CK(clk), .RN(n1569), .Q(
        \gbuff[17][28] ) );
  DFFRX1 \gbuff_reg[17][27]  ( .D(n2247), .CK(clk), .RN(n1569), .Q(
        \gbuff[17][27] ) );
  DFFRX1 \gbuff_reg[17][26]  ( .D(n2248), .CK(clk), .RN(n1569), .Q(
        \gbuff[17][26] ) );
  DFFRX1 \gbuff_reg[17][25]  ( .D(n2249), .CK(clk), .RN(n1569), .Q(
        \gbuff[17][25] ) );
  DFFRX1 \gbuff_reg[17][24]  ( .D(n2250), .CK(clk), .RN(n1569), .Q(
        \gbuff[17][24] ) );
  DFFRX1 \gbuff_reg[17][23]  ( .D(n2251), .CK(clk), .RN(n1569), .Q(
        \gbuff[17][23] ) );
  DFFRX1 \gbuff_reg[17][22]  ( .D(n2252), .CK(clk), .RN(n1569), .Q(
        \gbuff[17][22] ) );
  DFFRX1 \gbuff_reg[17][21]  ( .D(n2253), .CK(clk), .RN(n1569), .Q(
        \gbuff[17][21] ) );
  DFFRX1 \gbuff_reg[17][20]  ( .D(n2254), .CK(clk), .RN(n1569), .Q(
        \gbuff[17][20] ) );
  DFFRX1 \gbuff_reg[17][19]  ( .D(n2255), .CK(clk), .RN(n1568), .Q(
        \gbuff[17][19] ) );
  DFFRX1 \gbuff_reg[17][18]  ( .D(n2256), .CK(clk), .RN(n1568), .Q(
        \gbuff[17][18] ) );
  DFFRX1 \gbuff_reg[17][17]  ( .D(n2257), .CK(clk), .RN(n1568), .Q(
        \gbuff[17][17] ) );
  DFFRX1 \gbuff_reg[17][16]  ( .D(n2258), .CK(clk), .RN(n1568), .Q(
        \gbuff[17][16] ) );
  DFFRX1 \gbuff_reg[17][15]  ( .D(n2259), .CK(clk), .RN(n1568), .Q(
        \gbuff[17][15] ) );
  DFFRX1 \gbuff_reg[17][14]  ( .D(n2260), .CK(clk), .RN(n1568), .Q(
        \gbuff[17][14] ) );
  DFFRX1 \gbuff_reg[17][13]  ( .D(n2261), .CK(clk), .RN(n1568), .Q(
        \gbuff[17][13] ) );
  DFFRX1 \gbuff_reg[17][12]  ( .D(n2262), .CK(clk), .RN(n1568), .Q(
        \gbuff[17][12] ) );
  DFFRX1 \gbuff_reg[17][11]  ( .D(n2263), .CK(clk), .RN(n1568), .Q(
        \gbuff[17][11] ) );
  DFFRX1 \gbuff_reg[17][10]  ( .D(n2264), .CK(clk), .RN(n1568), .Q(
        \gbuff[17][10] ) );
  DFFRX1 \gbuff_reg[17][9]  ( .D(n2265), .CK(clk), .RN(n1568), .Q(
        \gbuff[17][9] ) );
  DFFRX1 \gbuff_reg[17][8]  ( .D(n2266), .CK(clk), .RN(n1568), .Q(
        \gbuff[17][8] ) );
  DFFRX1 \gbuff_reg[17][7]  ( .D(n2267), .CK(clk), .RN(n1567), .Q(
        \gbuff[17][7] ) );
  DFFRX1 \gbuff_reg[17][6]  ( .D(n2268), .CK(clk), .RN(n1567), .Q(
        \gbuff[17][6] ) );
  DFFRX1 \gbuff_reg[17][5]  ( .D(n2269), .CK(clk), .RN(n1567), .Q(
        \gbuff[17][5] ) );
  DFFRX1 \gbuff_reg[17][4]  ( .D(n2270), .CK(clk), .RN(n1567), .Q(
        \gbuff[17][4] ) );
  DFFRX1 \gbuff_reg[17][3]  ( .D(n2271), .CK(clk), .RN(n1567), .Q(
        \gbuff[17][3] ) );
  DFFRX1 \gbuff_reg[17][2]  ( .D(n2272), .CK(clk), .RN(n1567), .Q(
        \gbuff[17][2] ) );
  DFFRX1 \gbuff_reg[17][1]  ( .D(n2273), .CK(clk), .RN(n1567), .Q(
        \gbuff[17][1] ) );
  DFFRX1 \gbuff_reg[17][0]  ( .D(n2274), .CK(clk), .RN(n1567), .Q(
        \gbuff[17][0] ) );
  DFFRX1 \gbuff_reg[13][31]  ( .D(n2371), .CK(clk), .RN(n1559), .Q(
        \gbuff[13][31] ) );
  DFFRX1 \gbuff_reg[13][30]  ( .D(n2372), .CK(clk), .RN(n1559), .Q(
        \gbuff[13][30] ) );
  DFFRX1 \gbuff_reg[13][29]  ( .D(n2373), .CK(clk), .RN(n1559), .Q(
        \gbuff[13][29] ) );
  DFFRX1 \gbuff_reg[13][28]  ( .D(n2374), .CK(clk), .RN(n1559), .Q(
        \gbuff[13][28] ) );
  DFFRX1 \gbuff_reg[13][27]  ( .D(n2375), .CK(clk), .RN(n1558), .Q(
        \gbuff[13][27] ) );
  DFFRX1 \gbuff_reg[13][26]  ( .D(n2376), .CK(clk), .RN(n1558), .Q(
        \gbuff[13][26] ) );
  DFFRX1 \gbuff_reg[13][25]  ( .D(n2377), .CK(clk), .RN(n1558), .Q(
        \gbuff[13][25] ) );
  DFFRX1 \gbuff_reg[13][24]  ( .D(n2378), .CK(clk), .RN(n1558), .Q(
        \gbuff[13][24] ) );
  DFFRX1 \gbuff_reg[13][23]  ( .D(n2379), .CK(clk), .RN(n1558), .Q(
        \gbuff[13][23] ) );
  DFFRX1 \gbuff_reg[13][22]  ( .D(n2380), .CK(clk), .RN(n1558), .Q(
        \gbuff[13][22] ) );
  DFFRX1 \gbuff_reg[13][21]  ( .D(n2381), .CK(clk), .RN(n1558), .Q(
        \gbuff[13][21] ) );
  DFFRX1 \gbuff_reg[13][20]  ( .D(n2382), .CK(clk), .RN(n1558), .Q(
        \gbuff[13][20] ) );
  DFFRX1 \gbuff_reg[13][19]  ( .D(n2383), .CK(clk), .RN(n1558), .Q(
        \gbuff[13][19] ) );
  DFFRX1 \gbuff_reg[13][18]  ( .D(n2384), .CK(clk), .RN(n1558), .Q(
        \gbuff[13][18] ) );
  DFFRX1 \gbuff_reg[13][17]  ( .D(n2385), .CK(clk), .RN(n1558), .Q(
        \gbuff[13][17] ) );
  DFFRX1 \gbuff_reg[13][16]  ( .D(n2386), .CK(clk), .RN(n1558), .Q(
        \gbuff[13][16] ) );
  DFFRX1 \gbuff_reg[13][15]  ( .D(n2387), .CK(clk), .RN(n1557), .Q(
        \gbuff[13][15] ) );
  DFFRX1 \gbuff_reg[13][14]  ( .D(n2388), .CK(clk), .RN(n1557), .Q(
        \gbuff[13][14] ) );
  DFFRX1 \gbuff_reg[13][13]  ( .D(n2389), .CK(clk), .RN(n1557), .Q(
        \gbuff[13][13] ) );
  DFFRX1 \gbuff_reg[13][12]  ( .D(n2390), .CK(clk), .RN(n1557), .Q(
        \gbuff[13][12] ) );
  DFFRX1 \gbuff_reg[13][11]  ( .D(n2391), .CK(clk), .RN(n1557), .Q(
        \gbuff[13][11] ) );
  DFFRX1 \gbuff_reg[13][10]  ( .D(n2392), .CK(clk), .RN(n1557), .Q(
        \gbuff[13][10] ) );
  DFFRX1 \gbuff_reg[13][9]  ( .D(n2393), .CK(clk), .RN(n1557), .Q(
        \gbuff[13][9] ) );
  DFFRX1 \gbuff_reg[13][8]  ( .D(n2394), .CK(clk), .RN(n1557), .Q(
        \gbuff[13][8] ) );
  DFFRX1 \gbuff_reg[13][7]  ( .D(n2395), .CK(clk), .RN(n1557), .Q(
        \gbuff[13][7] ) );
  DFFRX1 \gbuff_reg[13][6]  ( .D(n2396), .CK(clk), .RN(n1557), .Q(
        \gbuff[13][6] ) );
  DFFRX1 \gbuff_reg[13][5]  ( .D(n2397), .CK(clk), .RN(n1557), .Q(
        \gbuff[13][5] ) );
  DFFRX1 \gbuff_reg[13][4]  ( .D(n2398), .CK(clk), .RN(n1557), .Q(
        \gbuff[13][4] ) );
  DFFRX1 \gbuff_reg[13][3]  ( .D(n2399), .CK(clk), .RN(n1556), .Q(
        \gbuff[13][3] ) );
  DFFRX1 \gbuff_reg[13][2]  ( .D(n2400), .CK(clk), .RN(n1556), .Q(
        \gbuff[13][2] ) );
  DFFRX1 \gbuff_reg[13][1]  ( .D(n2401), .CK(clk), .RN(n1556), .Q(
        \gbuff[13][1] ) );
  DFFRX1 \gbuff_reg[13][0]  ( .D(n2402), .CK(clk), .RN(n1556), .Q(
        \gbuff[13][0] ) );
  DFFRX1 \gbuff_reg[9][31]  ( .D(n2499), .CK(clk), .RN(n1548), .Q(
        \gbuff[9][31] ) );
  DFFRX1 \gbuff_reg[9][30]  ( .D(n2500), .CK(clk), .RN(n1548), .Q(
        \gbuff[9][30] ) );
  DFFRX1 \gbuff_reg[9][29]  ( .D(n2501), .CK(clk), .RN(n1548), .Q(
        \gbuff[9][29] ) );
  DFFRX1 \gbuff_reg[9][28]  ( .D(n2502), .CK(clk), .RN(n1548), .Q(
        \gbuff[9][28] ) );
  DFFRX1 \gbuff_reg[9][27]  ( .D(n2503), .CK(clk), .RN(n1548), .Q(
        \gbuff[9][27] ) );
  DFFRX1 \gbuff_reg[9][26]  ( .D(n2504), .CK(clk), .RN(n1548), .Q(
        \gbuff[9][26] ) );
  DFFRX1 \gbuff_reg[9][25]  ( .D(n2505), .CK(clk), .RN(n1548), .Q(
        \gbuff[9][25] ) );
  DFFRX1 \gbuff_reg[9][24]  ( .D(n2506), .CK(clk), .RN(n1548), .Q(
        \gbuff[9][24] ) );
  DFFRX1 \gbuff_reg[9][23]  ( .D(n2507), .CK(clk), .RN(n1547), .Q(
        \gbuff[9][23] ) );
  DFFRX1 \gbuff_reg[9][22]  ( .D(n2508), .CK(clk), .RN(n1547), .Q(
        \gbuff[9][22] ) );
  DFFRX1 \gbuff_reg[9][21]  ( .D(n2509), .CK(clk), .RN(n1547), .Q(
        \gbuff[9][21] ) );
  DFFRX1 \gbuff_reg[9][20]  ( .D(n2510), .CK(clk), .RN(n1547), .Q(
        \gbuff[9][20] ) );
  DFFRX1 \gbuff_reg[9][19]  ( .D(n2511), .CK(clk), .RN(n1547), .Q(
        \gbuff[9][19] ) );
  DFFRX1 \gbuff_reg[9][18]  ( .D(n2512), .CK(clk), .RN(n1547), .Q(
        \gbuff[9][18] ) );
  DFFRX1 \gbuff_reg[9][17]  ( .D(n2513), .CK(clk), .RN(n1547), .Q(
        \gbuff[9][17] ) );
  DFFRX1 \gbuff_reg[9][16]  ( .D(n2514), .CK(clk), .RN(n1547), .Q(
        \gbuff[9][16] ) );
  DFFRX1 \gbuff_reg[9][15]  ( .D(n2515), .CK(clk), .RN(n1547), .Q(
        \gbuff[9][15] ) );
  DFFRX1 \gbuff_reg[9][14]  ( .D(n2516), .CK(clk), .RN(n1547), .Q(
        \gbuff[9][14] ) );
  DFFRX1 \gbuff_reg[9][13]  ( .D(n2517), .CK(clk), .RN(n1547), .Q(
        \gbuff[9][13] ) );
  DFFRX1 \gbuff_reg[9][12]  ( .D(n2518), .CK(clk), .RN(n1547), .Q(
        \gbuff[9][12] ) );
  DFFRX1 \gbuff_reg[9][11]  ( .D(n2519), .CK(clk), .RN(n1546), .Q(
        \gbuff[9][11] ) );
  DFFRX1 \gbuff_reg[9][10]  ( .D(n2520), .CK(clk), .RN(n1546), .Q(
        \gbuff[9][10] ) );
  DFFRX1 \gbuff_reg[9][9]  ( .D(n2521), .CK(clk), .RN(n1546), .Q(\gbuff[9][9] ) );
  DFFRX1 \gbuff_reg[9][8]  ( .D(n2522), .CK(clk), .RN(n1546), .Q(\gbuff[9][8] ) );
  DFFRX1 \gbuff_reg[9][7]  ( .D(n2523), .CK(clk), .RN(n1546), .Q(\gbuff[9][7] ) );
  DFFRX1 \gbuff_reg[9][6]  ( .D(n2524), .CK(clk), .RN(n1546), .Q(\gbuff[9][6] ) );
  DFFRX1 \gbuff_reg[9][5]  ( .D(n2525), .CK(clk), .RN(n1546), .Q(\gbuff[9][5] ) );
  DFFRX1 \gbuff_reg[9][4]  ( .D(n2526), .CK(clk), .RN(n1546), .Q(\gbuff[9][4] ) );
  DFFRX1 \gbuff_reg[9][3]  ( .D(n2527), .CK(clk), .RN(n1546), .Q(\gbuff[9][3] ) );
  DFFRX1 \gbuff_reg[9][2]  ( .D(n2528), .CK(clk), .RN(n1546), .Q(\gbuff[9][2] ) );
  DFFRX1 \gbuff_reg[9][1]  ( .D(n2529), .CK(clk), .RN(n1546), .Q(\gbuff[9][1] ) );
  DFFRX1 \gbuff_reg[9][0]  ( .D(n2530), .CK(clk), .RN(n1546), .Q(\gbuff[9][0] ) );
  DFFRX1 \gbuff_reg[5][31]  ( .D(n2627), .CK(clk), .RN(n1537), .Q(
        \gbuff[5][31] ) );
  DFFRX1 \gbuff_reg[5][30]  ( .D(n2628), .CK(clk), .RN(n1537), .Q(
        \gbuff[5][30] ) );
  DFFRX1 \gbuff_reg[5][29]  ( .D(n2629), .CK(clk), .RN(n1537), .Q(
        \gbuff[5][29] ) );
  DFFRX1 \gbuff_reg[5][28]  ( .D(n2630), .CK(clk), .RN(n1537), .Q(
        \gbuff[5][28] ) );
  DFFRX1 \gbuff_reg[5][27]  ( .D(n2631), .CK(clk), .RN(n1537), .Q(
        \gbuff[5][27] ) );
  DFFRX1 \gbuff_reg[5][26]  ( .D(n2632), .CK(clk), .RN(n1537), .Q(
        \gbuff[5][26] ) );
  DFFRX1 \gbuff_reg[5][25]  ( .D(n2633), .CK(clk), .RN(n1537), .Q(
        \gbuff[5][25] ) );
  DFFRX1 \gbuff_reg[5][24]  ( .D(n2634), .CK(clk), .RN(n1537), .Q(
        \gbuff[5][24] ) );
  DFFRX1 \gbuff_reg[5][23]  ( .D(n2635), .CK(clk), .RN(n1537), .Q(
        \gbuff[5][23] ) );
  DFFRX1 \gbuff_reg[5][22]  ( .D(n2636), .CK(clk), .RN(n1537), .Q(
        \gbuff[5][22] ) );
  DFFRX1 \gbuff_reg[5][21]  ( .D(n2637), .CK(clk), .RN(n1537), .Q(
        \gbuff[5][21] ) );
  DFFRX1 \gbuff_reg[5][20]  ( .D(n2638), .CK(clk), .RN(n1537), .Q(
        \gbuff[5][20] ) );
  DFFRX1 \gbuff_reg[5][19]  ( .D(n2639), .CK(clk), .RN(n1536), .Q(
        \gbuff[5][19] ) );
  DFFRX1 \gbuff_reg[5][18]  ( .D(n2640), .CK(clk), .RN(n1536), .Q(
        \gbuff[5][18] ) );
  DFFRX1 \gbuff_reg[5][17]  ( .D(n2641), .CK(clk), .RN(n1536), .Q(
        \gbuff[5][17] ) );
  DFFRX1 \gbuff_reg[5][16]  ( .D(n2642), .CK(clk), .RN(n1536), .Q(
        \gbuff[5][16] ) );
  DFFRX1 \gbuff_reg[5][15]  ( .D(n2643), .CK(clk), .RN(n1536), .Q(
        \gbuff[5][15] ) );
  DFFRX1 \gbuff_reg[5][14]  ( .D(n2644), .CK(clk), .RN(n1536), .Q(
        \gbuff[5][14] ) );
  DFFRX1 \gbuff_reg[5][13]  ( .D(n2645), .CK(clk), .RN(n1536), .Q(
        \gbuff[5][13] ) );
  DFFRX1 \gbuff_reg[5][12]  ( .D(n2646), .CK(clk), .RN(n1536), .Q(
        \gbuff[5][12] ) );
  DFFRX1 \gbuff_reg[5][11]  ( .D(n2647), .CK(clk), .RN(n1536), .Q(
        \gbuff[5][11] ) );
  DFFRX1 \gbuff_reg[5][10]  ( .D(n2648), .CK(clk), .RN(n1536), .Q(
        \gbuff[5][10] ) );
  DFFRX1 \gbuff_reg[5][9]  ( .D(n2649), .CK(clk), .RN(n1536), .Q(\gbuff[5][9] ) );
  DFFRX1 \gbuff_reg[5][8]  ( .D(n2650), .CK(clk), .RN(n1536), .Q(\gbuff[5][8] ) );
  DFFRX1 \gbuff_reg[5][7]  ( .D(n2651), .CK(clk), .RN(n1535), .Q(\gbuff[5][7] ) );
  DFFRX1 \gbuff_reg[5][6]  ( .D(n2652), .CK(clk), .RN(n1535), .Q(\gbuff[5][6] ) );
  DFFRX1 \gbuff_reg[5][5]  ( .D(n2653), .CK(clk), .RN(n1535), .Q(\gbuff[5][5] ) );
  DFFRX1 \gbuff_reg[5][4]  ( .D(n2654), .CK(clk), .RN(n1535), .Q(\gbuff[5][4] ) );
  DFFRX1 \gbuff_reg[5][3]  ( .D(n2655), .CK(clk), .RN(n1535), .Q(\gbuff[5][3] ) );
  DFFRX1 \gbuff_reg[5][2]  ( .D(n2656), .CK(clk), .RN(n1535), .Q(\gbuff[5][2] ) );
  DFFRX1 \gbuff_reg[5][1]  ( .D(n2657), .CK(clk), .RN(n1535), .Q(\gbuff[5][1] ) );
  DFFRX1 \gbuff_reg[5][0]  ( .D(n2658), .CK(clk), .RN(n1535), .Q(\gbuff[5][0] ) );
  DFFRX1 \gbuff_reg[1][31]  ( .D(n2755), .CK(clk), .RN(n1527), .Q(
        \gbuff[1][31] ) );
  DFFRX1 \gbuff_reg[1][30]  ( .D(n2756), .CK(clk), .RN(n1527), .Q(
        \gbuff[1][30] ) );
  DFFRX1 \gbuff_reg[1][29]  ( .D(n2757), .CK(clk), .RN(n1527), .Q(
        \gbuff[1][29] ) );
  DFFRX1 \gbuff_reg[1][28]  ( .D(n2758), .CK(clk), .RN(n1527), .Q(
        \gbuff[1][28] ) );
  DFFRX1 \gbuff_reg[1][27]  ( .D(n2759), .CK(clk), .RN(n1526), .Q(
        \gbuff[1][27] ) );
  DFFRX1 \gbuff_reg[1][26]  ( .D(n2760), .CK(clk), .RN(n1526), .Q(
        \gbuff[1][26] ) );
  DFFRX1 \gbuff_reg[1][25]  ( .D(n2761), .CK(clk), .RN(n1526), .Q(
        \gbuff[1][25] ) );
  DFFRX1 \gbuff_reg[1][24]  ( .D(n2762), .CK(clk), .RN(n1526), .Q(
        \gbuff[1][24] ) );
  DFFRX1 \gbuff_reg[1][23]  ( .D(n2763), .CK(clk), .RN(n1526), .Q(
        \gbuff[1][23] ) );
  DFFRX1 \gbuff_reg[1][22]  ( .D(n2764), .CK(clk), .RN(n1526), .Q(
        \gbuff[1][22] ) );
  DFFRX1 \gbuff_reg[1][21]  ( .D(n2765), .CK(clk), .RN(n1526), .Q(
        \gbuff[1][21] ) );
  DFFRX1 \gbuff_reg[1][20]  ( .D(n2766), .CK(clk), .RN(n1526), .Q(
        \gbuff[1][20] ) );
  DFFRX1 \gbuff_reg[1][19]  ( .D(n2767), .CK(clk), .RN(n1526), .Q(
        \gbuff[1][19] ) );
  DFFRX1 \gbuff_reg[1][18]  ( .D(n2768), .CK(clk), .RN(n1526), .Q(
        \gbuff[1][18] ) );
  DFFRX1 \gbuff_reg[1][17]  ( .D(n2769), .CK(clk), .RN(n1526), .Q(
        \gbuff[1][17] ) );
  DFFRX1 \gbuff_reg[1][16]  ( .D(n2770), .CK(clk), .RN(n1526), .Q(
        \gbuff[1][16] ) );
  DFFRX1 \gbuff_reg[1][15]  ( .D(n2771), .CK(clk), .RN(n1525), .Q(
        \gbuff[1][15] ) );
  DFFRX1 \gbuff_reg[1][14]  ( .D(n2772), .CK(clk), .RN(n1525), .Q(
        \gbuff[1][14] ) );
  DFFRX1 \gbuff_reg[1][13]  ( .D(n2773), .CK(clk), .RN(n1525), .Q(
        \gbuff[1][13] ) );
  DFFRX1 \gbuff_reg[1][12]  ( .D(n2774), .CK(clk), .RN(n1525), .Q(
        \gbuff[1][12] ) );
  DFFRX1 \gbuff_reg[1][11]  ( .D(n2775), .CK(clk), .RN(n1525), .Q(
        \gbuff[1][11] ) );
  DFFRX1 \gbuff_reg[1][10]  ( .D(n2776), .CK(clk), .RN(n1525), .Q(
        \gbuff[1][10] ) );
  DFFRX1 \gbuff_reg[1][9]  ( .D(n2777), .CK(clk), .RN(n1525), .Q(\gbuff[1][9] ) );
  DFFRX1 \gbuff_reg[1][8]  ( .D(n2778), .CK(clk), .RN(n1525), .Q(\gbuff[1][8] ) );
  DFFRX1 \gbuff_reg[1][7]  ( .D(n2779), .CK(clk), .RN(n1525), .Q(\gbuff[1][7] ) );
  DFFRX1 \gbuff_reg[1][6]  ( .D(n2780), .CK(clk), .RN(n1525), .Q(\gbuff[1][6] ) );
  DFFRX1 \gbuff_reg[1][5]  ( .D(n2781), .CK(clk), .RN(n1525), .Q(\gbuff[1][5] ) );
  DFFRX1 \gbuff_reg[1][4]  ( .D(n2782), .CK(clk), .RN(n1525), .Q(\gbuff[1][4] ) );
  DFFRX1 \gbuff_reg[1][3]  ( .D(n2783), .CK(clk), .RN(n1524), .Q(\gbuff[1][3] ) );
  DFFRX1 \gbuff_reg[1][2]  ( .D(n2784), .CK(clk), .RN(n1524), .Q(\gbuff[1][2] ) );
  DFFRX1 \gbuff_reg[1][1]  ( .D(n2785), .CK(clk), .RN(n1524), .Q(\gbuff[1][1] ) );
  DFFRX1 \gbuff_reg[1][0]  ( .D(n2786), .CK(clk), .RN(n1524), .Q(\gbuff[1][0] ) );
  DFFRX1 \gbuff_reg[31][31]  ( .D(n1795), .CK(clk), .RN(n1607), .Q(
        \gbuff[31][31] ) );
  DFFRX1 \gbuff_reg[31][30]  ( .D(n1796), .CK(clk), .RN(n1607), .Q(
        \gbuff[31][30] ) );
  DFFRX1 \gbuff_reg[31][29]  ( .D(n1797), .CK(clk), .RN(n1607), .Q(
        \gbuff[31][29] ) );
  DFFRX1 \gbuff_reg[31][28]  ( .D(n1798), .CK(clk), .RN(n1607), .Q(
        \gbuff[31][28] ) );
  DFFRX1 \gbuff_reg[31][27]  ( .D(n1799), .CK(clk), .RN(n1606), .Q(
        \gbuff[31][27] ) );
  DFFRX1 \gbuff_reg[31][26]  ( .D(n1800), .CK(clk), .RN(n1606), .Q(
        \gbuff[31][26] ) );
  DFFRX1 \gbuff_reg[31][25]  ( .D(n1801), .CK(clk), .RN(n1606), .Q(
        \gbuff[31][25] ) );
  DFFRX1 \gbuff_reg[31][24]  ( .D(n1802), .CK(clk), .RN(n1606), .Q(
        \gbuff[31][24] ) );
  DFFRX1 \gbuff_reg[31][23]  ( .D(n1803), .CK(clk), .RN(n1606), .Q(
        \gbuff[31][23] ) );
  DFFRX1 \gbuff_reg[31][22]  ( .D(n1804), .CK(clk), .RN(n1606), .Q(
        \gbuff[31][22] ) );
  DFFRX1 \gbuff_reg[31][21]  ( .D(n1805), .CK(clk), .RN(n1606), .Q(
        \gbuff[31][21] ) );
  DFFRX1 \gbuff_reg[31][20]  ( .D(n1806), .CK(clk), .RN(n1606), .Q(
        \gbuff[31][20] ) );
  DFFRX1 \gbuff_reg[31][19]  ( .D(n1807), .CK(clk), .RN(n1606), .Q(
        \gbuff[31][19] ) );
  DFFRX1 \gbuff_reg[31][18]  ( .D(n1808), .CK(clk), .RN(n1606), .Q(
        \gbuff[31][18] ) );
  DFFRX1 \gbuff_reg[31][17]  ( .D(n1809), .CK(clk), .RN(n1606), .Q(
        \gbuff[31][17] ) );
  DFFRX1 \gbuff_reg[31][16]  ( .D(n1810), .CK(clk), .RN(n1606), .Q(
        \gbuff[31][16] ) );
  DFFRX1 \gbuff_reg[31][15]  ( .D(n1811), .CK(clk), .RN(n1605), .Q(
        \gbuff[31][15] ) );
  DFFRX1 \gbuff_reg[31][14]  ( .D(n1812), .CK(clk), .RN(n1605), .Q(
        \gbuff[31][14] ) );
  DFFRX1 \gbuff_reg[31][13]  ( .D(n1813), .CK(clk), .RN(n1605), .Q(
        \gbuff[31][13] ) );
  DFFRX1 \gbuff_reg[31][12]  ( .D(n1814), .CK(clk), .RN(n1605), .Q(
        \gbuff[31][12] ) );
  DFFRX1 \gbuff_reg[31][11]  ( .D(n1815), .CK(clk), .RN(n1605), .Q(
        \gbuff[31][11] ) );
  DFFRX1 \gbuff_reg[31][10]  ( .D(n1816), .CK(clk), .RN(n1605), .Q(
        \gbuff[31][10] ) );
  DFFRX1 \gbuff_reg[31][9]  ( .D(n1817), .CK(clk), .RN(n1605), .Q(
        \gbuff[31][9] ) );
  DFFRX1 \gbuff_reg[31][8]  ( .D(n1818), .CK(clk), .RN(n1605), .Q(
        \gbuff[31][8] ) );
  DFFRX1 \gbuff_reg[31][7]  ( .D(n1819), .CK(clk), .RN(n1605), .Q(
        \gbuff[31][7] ) );
  DFFRX1 \gbuff_reg[31][6]  ( .D(n1820), .CK(clk), .RN(n1605), .Q(
        \gbuff[31][6] ) );
  DFFRX1 \gbuff_reg[31][5]  ( .D(n1821), .CK(clk), .RN(n1605), .Q(
        \gbuff[31][5] ) );
  DFFRX1 \gbuff_reg[31][4]  ( .D(n1822), .CK(clk), .RN(n1605), .Q(
        \gbuff[31][4] ) );
  DFFRX1 \gbuff_reg[31][3]  ( .D(n1823), .CK(clk), .RN(n1604), .Q(
        \gbuff[31][3] ) );
  DFFRX1 \gbuff_reg[31][2]  ( .D(n1824), .CK(clk), .RN(n1604), .Q(
        \gbuff[31][2] ) );
  DFFRX1 \gbuff_reg[31][1]  ( .D(n1825), .CK(clk), .RN(n1604), .Q(
        \gbuff[31][1] ) );
  DFFRX1 \gbuff_reg[31][0]  ( .D(n1826), .CK(clk), .RN(n1604), .Q(
        \gbuff[31][0] ) );
  DFFRX1 \gbuff_reg[27][31]  ( .D(n1923), .CK(clk), .RN(n1596), .Q(
        \gbuff[27][31] ) );
  DFFRX1 \gbuff_reg[27][30]  ( .D(n1924), .CK(clk), .RN(n1596), .Q(
        \gbuff[27][30] ) );
  DFFRX1 \gbuff_reg[27][29]  ( .D(n1925), .CK(clk), .RN(n1596), .Q(
        \gbuff[27][29] ) );
  DFFRX1 \gbuff_reg[27][28]  ( .D(n1926), .CK(clk), .RN(n1596), .Q(
        \gbuff[27][28] ) );
  DFFRX1 \gbuff_reg[27][27]  ( .D(n1927), .CK(clk), .RN(n1596), .Q(
        \gbuff[27][27] ) );
  DFFRX1 \gbuff_reg[27][26]  ( .D(n1928), .CK(clk), .RN(n1596), .Q(
        \gbuff[27][26] ) );
  DFFRX1 \gbuff_reg[27][25]  ( .D(n1929), .CK(clk), .RN(n1596), .Q(
        \gbuff[27][25] ) );
  DFFRX1 \gbuff_reg[27][24]  ( .D(n1930), .CK(clk), .RN(n1596), .Q(
        \gbuff[27][24] ) );
  DFFRX1 \gbuff_reg[27][23]  ( .D(n1931), .CK(clk), .RN(n1595), .Q(
        \gbuff[27][23] ) );
  DFFRX1 \gbuff_reg[27][22]  ( .D(n1932), .CK(clk), .RN(n1595), .Q(
        \gbuff[27][22] ) );
  DFFRX1 \gbuff_reg[27][21]  ( .D(n1933), .CK(clk), .RN(n1595), .Q(
        \gbuff[27][21] ) );
  DFFRX1 \gbuff_reg[27][20]  ( .D(n1934), .CK(clk), .RN(n1595), .Q(
        \gbuff[27][20] ) );
  DFFRX1 \gbuff_reg[27][19]  ( .D(n1935), .CK(clk), .RN(n1595), .Q(
        \gbuff[27][19] ) );
  DFFRX1 \gbuff_reg[27][18]  ( .D(n1936), .CK(clk), .RN(n1595), .Q(
        \gbuff[27][18] ) );
  DFFRX1 \gbuff_reg[27][17]  ( .D(n1937), .CK(clk), .RN(n1595), .Q(
        \gbuff[27][17] ) );
  DFFRX1 \gbuff_reg[27][16]  ( .D(n1938), .CK(clk), .RN(n1595), .Q(
        \gbuff[27][16] ) );
  DFFRX1 \gbuff_reg[27][15]  ( .D(n1939), .CK(clk), .RN(n1595), .Q(
        \gbuff[27][15] ) );
  DFFRX1 \gbuff_reg[27][14]  ( .D(n1940), .CK(clk), .RN(n1595), .Q(
        \gbuff[27][14] ) );
  DFFRX1 \gbuff_reg[27][13]  ( .D(n1941), .CK(clk), .RN(n1595), .Q(
        \gbuff[27][13] ) );
  DFFRX1 \gbuff_reg[27][12]  ( .D(n1942), .CK(clk), .RN(n1595), .Q(
        \gbuff[27][12] ) );
  DFFRX1 \gbuff_reg[27][11]  ( .D(n1943), .CK(clk), .RN(n1594), .Q(
        \gbuff[27][11] ) );
  DFFRX1 \gbuff_reg[27][10]  ( .D(n1944), .CK(clk), .RN(n1594), .Q(
        \gbuff[27][10] ) );
  DFFRX1 \gbuff_reg[27][9]  ( .D(n1945), .CK(clk), .RN(n1594), .Q(
        \gbuff[27][9] ) );
  DFFRX1 \gbuff_reg[27][8]  ( .D(n1946), .CK(clk), .RN(n1594), .Q(
        \gbuff[27][8] ) );
  DFFRX1 \gbuff_reg[27][7]  ( .D(n1947), .CK(clk), .RN(n1594), .Q(
        \gbuff[27][7] ) );
  DFFRX1 \gbuff_reg[27][6]  ( .D(n1948), .CK(clk), .RN(n1594), .Q(
        \gbuff[27][6] ) );
  DFFRX1 \gbuff_reg[27][5]  ( .D(n1949), .CK(clk), .RN(n1594), .Q(
        \gbuff[27][5] ) );
  DFFRX1 \gbuff_reg[27][4]  ( .D(n1950), .CK(clk), .RN(n1594), .Q(
        \gbuff[27][4] ) );
  DFFRX1 \gbuff_reg[27][3]  ( .D(n1951), .CK(clk), .RN(n1594), .Q(
        \gbuff[27][3] ) );
  DFFRX1 \gbuff_reg[27][2]  ( .D(n1952), .CK(clk), .RN(n1594), .Q(
        \gbuff[27][2] ) );
  DFFRX1 \gbuff_reg[27][1]  ( .D(n1953), .CK(clk), .RN(n1594), .Q(
        \gbuff[27][1] ) );
  DFFRX1 \gbuff_reg[27][0]  ( .D(n1954), .CK(clk), .RN(n1594), .Q(
        \gbuff[27][0] ) );
  DFFRX1 \gbuff_reg[23][31]  ( .D(n2051), .CK(clk), .RN(n1585), .Q(
        \gbuff[23][31] ) );
  DFFRX1 \gbuff_reg[23][30]  ( .D(n2052), .CK(clk), .RN(n1585), .Q(
        \gbuff[23][30] ) );
  DFFRX1 \gbuff_reg[23][29]  ( .D(n2053), .CK(clk), .RN(n1585), .Q(
        \gbuff[23][29] ) );
  DFFRX1 \gbuff_reg[23][28]  ( .D(n2054), .CK(clk), .RN(n1585), .Q(
        \gbuff[23][28] ) );
  DFFRX1 \gbuff_reg[23][27]  ( .D(n2055), .CK(clk), .RN(n1585), .Q(
        \gbuff[23][27] ) );
  DFFRX1 \gbuff_reg[23][26]  ( .D(n2056), .CK(clk), .RN(n1585), .Q(
        \gbuff[23][26] ) );
  DFFRX1 \gbuff_reg[23][25]  ( .D(n2057), .CK(clk), .RN(n1585), .Q(
        \gbuff[23][25] ) );
  DFFRX1 \gbuff_reg[23][24]  ( .D(n2058), .CK(clk), .RN(n1585), .Q(
        \gbuff[23][24] ) );
  DFFRX1 \gbuff_reg[23][23]  ( .D(n2059), .CK(clk), .RN(n1585), .Q(
        \gbuff[23][23] ) );
  DFFRX1 \gbuff_reg[23][22]  ( .D(n2060), .CK(clk), .RN(n1585), .Q(
        \gbuff[23][22] ) );
  DFFRX1 \gbuff_reg[23][21]  ( .D(n2061), .CK(clk), .RN(n1585), .Q(
        \gbuff[23][21] ) );
  DFFRX1 \gbuff_reg[23][20]  ( .D(n2062), .CK(clk), .RN(n1585), .Q(
        \gbuff[23][20] ) );
  DFFRX1 \gbuff_reg[23][19]  ( .D(n2063), .CK(clk), .RN(n1584), .Q(
        \gbuff[23][19] ) );
  DFFRX1 \gbuff_reg[23][18]  ( .D(n2064), .CK(clk), .RN(n1584), .Q(
        \gbuff[23][18] ) );
  DFFRX1 \gbuff_reg[23][17]  ( .D(n2065), .CK(clk), .RN(n1584), .Q(
        \gbuff[23][17] ) );
  DFFRX1 \gbuff_reg[23][16]  ( .D(n2066), .CK(clk), .RN(n1584), .Q(
        \gbuff[23][16] ) );
  DFFRX1 \gbuff_reg[23][15]  ( .D(n2067), .CK(clk), .RN(n1584), .Q(
        \gbuff[23][15] ) );
  DFFRX1 \gbuff_reg[23][14]  ( .D(n2068), .CK(clk), .RN(n1584), .Q(
        \gbuff[23][14] ) );
  DFFRX1 \gbuff_reg[23][13]  ( .D(n2069), .CK(clk), .RN(n1584), .Q(
        \gbuff[23][13] ) );
  DFFRX1 \gbuff_reg[23][12]  ( .D(n2070), .CK(clk), .RN(n1584), .Q(
        \gbuff[23][12] ) );
  DFFRX1 \gbuff_reg[23][11]  ( .D(n2071), .CK(clk), .RN(n1584), .Q(
        \gbuff[23][11] ) );
  DFFRX1 \gbuff_reg[23][10]  ( .D(n2072), .CK(clk), .RN(n1584), .Q(
        \gbuff[23][10] ) );
  DFFRX1 \gbuff_reg[23][9]  ( .D(n2073), .CK(clk), .RN(n1584), .Q(
        \gbuff[23][9] ) );
  DFFRX1 \gbuff_reg[23][8]  ( .D(n2074), .CK(clk), .RN(n1584), .Q(
        \gbuff[23][8] ) );
  DFFRX1 \gbuff_reg[23][7]  ( .D(n2075), .CK(clk), .RN(n1583), .Q(
        \gbuff[23][7] ) );
  DFFRX1 \gbuff_reg[23][6]  ( .D(n2076), .CK(clk), .RN(n1583), .Q(
        \gbuff[23][6] ) );
  DFFRX1 \gbuff_reg[23][5]  ( .D(n2077), .CK(clk), .RN(n1583), .Q(
        \gbuff[23][5] ) );
  DFFRX1 \gbuff_reg[23][4]  ( .D(n2078), .CK(clk), .RN(n1583), .Q(
        \gbuff[23][4] ) );
  DFFRX1 \gbuff_reg[23][3]  ( .D(n2079), .CK(clk), .RN(n1583), .Q(
        \gbuff[23][3] ) );
  DFFRX1 \gbuff_reg[23][2]  ( .D(n2080), .CK(clk), .RN(n1583), .Q(
        \gbuff[23][2] ) );
  DFFRX1 \gbuff_reg[23][1]  ( .D(n2081), .CK(clk), .RN(n1583), .Q(
        \gbuff[23][1] ) );
  DFFRX1 \gbuff_reg[23][0]  ( .D(n2082), .CK(clk), .RN(n1583), .Q(
        \gbuff[23][0] ) );
  DFFRX1 \gbuff_reg[19][31]  ( .D(n2179), .CK(clk), .RN(n1575), .Q(
        \gbuff[19][31] ) );
  DFFRX1 \gbuff_reg[19][30]  ( .D(n2180), .CK(clk), .RN(n1575), .Q(
        \gbuff[19][30] ) );
  DFFRX1 \gbuff_reg[19][29]  ( .D(n2181), .CK(clk), .RN(n1575), .Q(
        \gbuff[19][29] ) );
  DFFRX1 \gbuff_reg[19][28]  ( .D(n2182), .CK(clk), .RN(n1575), .Q(
        \gbuff[19][28] ) );
  DFFRX1 \gbuff_reg[19][27]  ( .D(n2183), .CK(clk), .RN(n1574), .Q(
        \gbuff[19][27] ) );
  DFFRX1 \gbuff_reg[19][26]  ( .D(n2184), .CK(clk), .RN(n1574), .Q(
        \gbuff[19][26] ) );
  DFFRX1 \gbuff_reg[19][25]  ( .D(n2185), .CK(clk), .RN(n1574), .Q(
        \gbuff[19][25] ) );
  DFFRX1 \gbuff_reg[19][24]  ( .D(n2186), .CK(clk), .RN(n1574), .Q(
        \gbuff[19][24] ) );
  DFFRX1 \gbuff_reg[19][23]  ( .D(n2187), .CK(clk), .RN(n1574), .Q(
        \gbuff[19][23] ) );
  DFFRX1 \gbuff_reg[19][22]  ( .D(n2188), .CK(clk), .RN(n1574), .Q(
        \gbuff[19][22] ) );
  DFFRX1 \gbuff_reg[19][21]  ( .D(n2189), .CK(clk), .RN(n1574), .Q(
        \gbuff[19][21] ) );
  DFFRX1 \gbuff_reg[19][20]  ( .D(n2190), .CK(clk), .RN(n1574), .Q(
        \gbuff[19][20] ) );
  DFFRX1 \gbuff_reg[19][19]  ( .D(n2191), .CK(clk), .RN(n1574), .Q(
        \gbuff[19][19] ) );
  DFFRX1 \gbuff_reg[19][18]  ( .D(n2192), .CK(clk), .RN(n1574), .Q(
        \gbuff[19][18] ) );
  DFFRX1 \gbuff_reg[19][17]  ( .D(n2193), .CK(clk), .RN(n1574), .Q(
        \gbuff[19][17] ) );
  DFFRX1 \gbuff_reg[19][16]  ( .D(n2194), .CK(clk), .RN(n1574), .Q(
        \gbuff[19][16] ) );
  DFFRX1 \gbuff_reg[19][15]  ( .D(n2195), .CK(clk), .RN(n1573), .Q(
        \gbuff[19][15] ) );
  DFFRX1 \gbuff_reg[19][14]  ( .D(n2196), .CK(clk), .RN(n1573), .Q(
        \gbuff[19][14] ) );
  DFFRX1 \gbuff_reg[19][13]  ( .D(n2197), .CK(clk), .RN(n1573), .Q(
        \gbuff[19][13] ) );
  DFFRX1 \gbuff_reg[19][12]  ( .D(n2198), .CK(clk), .RN(n1573), .Q(
        \gbuff[19][12] ) );
  DFFRX1 \gbuff_reg[19][11]  ( .D(n2199), .CK(clk), .RN(n1573), .Q(
        \gbuff[19][11] ) );
  DFFRX1 \gbuff_reg[19][10]  ( .D(n2200), .CK(clk), .RN(n1573), .Q(
        \gbuff[19][10] ) );
  DFFRX1 \gbuff_reg[19][9]  ( .D(n2201), .CK(clk), .RN(n1573), .Q(
        \gbuff[19][9] ) );
  DFFRX1 \gbuff_reg[19][8]  ( .D(n2202), .CK(clk), .RN(n1573), .Q(
        \gbuff[19][8] ) );
  DFFRX1 \gbuff_reg[19][7]  ( .D(n2203), .CK(clk), .RN(n1573), .Q(
        \gbuff[19][7] ) );
  DFFRX1 \gbuff_reg[19][6]  ( .D(n2204), .CK(clk), .RN(n1573), .Q(
        \gbuff[19][6] ) );
  DFFRX1 \gbuff_reg[19][5]  ( .D(n2205), .CK(clk), .RN(n1573), .Q(
        \gbuff[19][5] ) );
  DFFRX1 \gbuff_reg[19][4]  ( .D(n2206), .CK(clk), .RN(n1573), .Q(
        \gbuff[19][4] ) );
  DFFRX1 \gbuff_reg[19][3]  ( .D(n2207), .CK(clk), .RN(n1572), .Q(
        \gbuff[19][3] ) );
  DFFRX1 \gbuff_reg[19][2]  ( .D(n2208), .CK(clk), .RN(n1572), .Q(
        \gbuff[19][2] ) );
  DFFRX1 \gbuff_reg[19][1]  ( .D(n2209), .CK(clk), .RN(n1572), .Q(
        \gbuff[19][1] ) );
  DFFRX1 \gbuff_reg[19][0]  ( .D(n2210), .CK(clk), .RN(n1572), .Q(
        \gbuff[19][0] ) );
  DFFRX1 \gbuff_reg[15][31]  ( .D(n2307), .CK(clk), .RN(n1564), .Q(
        \gbuff[15][31] ) );
  DFFRX1 \gbuff_reg[15][30]  ( .D(n2308), .CK(clk), .RN(n1564), .Q(
        \gbuff[15][30] ) );
  DFFRX1 \gbuff_reg[15][29]  ( .D(n2309), .CK(clk), .RN(n1564), .Q(
        \gbuff[15][29] ) );
  DFFRX1 \gbuff_reg[15][28]  ( .D(n2310), .CK(clk), .RN(n1564), .Q(
        \gbuff[15][28] ) );
  DFFRX1 \gbuff_reg[15][27]  ( .D(n2311), .CK(clk), .RN(n1564), .Q(
        \gbuff[15][27] ) );
  DFFRX1 \gbuff_reg[15][26]  ( .D(n2312), .CK(clk), .RN(n1564), .Q(
        \gbuff[15][26] ) );
  DFFRX1 \gbuff_reg[15][25]  ( .D(n2313), .CK(clk), .RN(n1564), .Q(
        \gbuff[15][25] ) );
  DFFRX1 \gbuff_reg[15][24]  ( .D(n2314), .CK(clk), .RN(n1564), .Q(
        \gbuff[15][24] ) );
  DFFRX1 \gbuff_reg[15][23]  ( .D(n2315), .CK(clk), .RN(n1563), .Q(
        \gbuff[15][23] ) );
  DFFRX1 \gbuff_reg[15][22]  ( .D(n2316), .CK(clk), .RN(n1563), .Q(
        \gbuff[15][22] ) );
  DFFRX1 \gbuff_reg[15][21]  ( .D(n2317), .CK(clk), .RN(n1563), .Q(
        \gbuff[15][21] ) );
  DFFRX1 \gbuff_reg[15][20]  ( .D(n2318), .CK(clk), .RN(n1563), .Q(
        \gbuff[15][20] ) );
  DFFRX1 \gbuff_reg[15][19]  ( .D(n2319), .CK(clk), .RN(n1563), .Q(
        \gbuff[15][19] ) );
  DFFRX1 \gbuff_reg[15][18]  ( .D(n2320), .CK(clk), .RN(n1563), .Q(
        \gbuff[15][18] ) );
  DFFRX1 \gbuff_reg[15][17]  ( .D(n2321), .CK(clk), .RN(n1563), .Q(
        \gbuff[15][17] ) );
  DFFRX1 \gbuff_reg[15][16]  ( .D(n2322), .CK(clk), .RN(n1563), .Q(
        \gbuff[15][16] ) );
  DFFRX1 \gbuff_reg[15][15]  ( .D(n2323), .CK(clk), .RN(n1563), .Q(
        \gbuff[15][15] ) );
  DFFRX1 \gbuff_reg[15][14]  ( .D(n2324), .CK(clk), .RN(n1563), .Q(
        \gbuff[15][14] ) );
  DFFRX1 \gbuff_reg[15][13]  ( .D(n2325), .CK(clk), .RN(n1563), .Q(
        \gbuff[15][13] ) );
  DFFRX1 \gbuff_reg[15][12]  ( .D(n2326), .CK(clk), .RN(n1563), .Q(
        \gbuff[15][12] ) );
  DFFRX1 \gbuff_reg[15][11]  ( .D(n2327), .CK(clk), .RN(n1562), .Q(
        \gbuff[15][11] ) );
  DFFRX1 \gbuff_reg[15][10]  ( .D(n2328), .CK(clk), .RN(n1562), .Q(
        \gbuff[15][10] ) );
  DFFRX1 \gbuff_reg[15][9]  ( .D(n2329), .CK(clk), .RN(n1562), .Q(
        \gbuff[15][9] ) );
  DFFRX1 \gbuff_reg[15][8]  ( .D(n2330), .CK(clk), .RN(n1562), .Q(
        \gbuff[15][8] ) );
  DFFRX1 \gbuff_reg[15][7]  ( .D(n2331), .CK(clk), .RN(n1562), .Q(
        \gbuff[15][7] ) );
  DFFRX1 \gbuff_reg[15][6]  ( .D(n2332), .CK(clk), .RN(n1562), .Q(
        \gbuff[15][6] ) );
  DFFRX1 \gbuff_reg[15][5]  ( .D(n2333), .CK(clk), .RN(n1562), .Q(
        \gbuff[15][5] ) );
  DFFRX1 \gbuff_reg[15][4]  ( .D(n2334), .CK(clk), .RN(n1562), .Q(
        \gbuff[15][4] ) );
  DFFRX1 \gbuff_reg[15][3]  ( .D(n2335), .CK(clk), .RN(n1562), .Q(
        \gbuff[15][3] ) );
  DFFRX1 \gbuff_reg[15][2]  ( .D(n2336), .CK(clk), .RN(n1562), .Q(
        \gbuff[15][2] ) );
  DFFRX1 \gbuff_reg[15][1]  ( .D(n2337), .CK(clk), .RN(n1562), .Q(
        \gbuff[15][1] ) );
  DFFRX1 \gbuff_reg[15][0]  ( .D(n2338), .CK(clk), .RN(n1562), .Q(
        \gbuff[15][0] ) );
  DFFRX1 \gbuff_reg[11][31]  ( .D(n2435), .CK(clk), .RN(n1553), .Q(
        \gbuff[11][31] ) );
  DFFRX1 \gbuff_reg[11][30]  ( .D(n2436), .CK(clk), .RN(n1553), .Q(
        \gbuff[11][30] ) );
  DFFRX1 \gbuff_reg[11][29]  ( .D(n2437), .CK(clk), .RN(n1553), .Q(
        \gbuff[11][29] ) );
  DFFRX1 \gbuff_reg[11][28]  ( .D(n2438), .CK(clk), .RN(n1553), .Q(
        \gbuff[11][28] ) );
  DFFRX1 \gbuff_reg[11][27]  ( .D(n2439), .CK(clk), .RN(n1553), .Q(
        \gbuff[11][27] ) );
  DFFRX1 \gbuff_reg[11][26]  ( .D(n2440), .CK(clk), .RN(n1553), .Q(
        \gbuff[11][26] ) );
  DFFRX1 \gbuff_reg[11][25]  ( .D(n2441), .CK(clk), .RN(n1553), .Q(
        \gbuff[11][25] ) );
  DFFRX1 \gbuff_reg[11][24]  ( .D(n2442), .CK(clk), .RN(n1553), .Q(
        \gbuff[11][24] ) );
  DFFRX1 \gbuff_reg[11][23]  ( .D(n2443), .CK(clk), .RN(n1553), .Q(
        \gbuff[11][23] ) );
  DFFRX1 \gbuff_reg[11][22]  ( .D(n2444), .CK(clk), .RN(n1553), .Q(
        \gbuff[11][22] ) );
  DFFRX1 \gbuff_reg[11][21]  ( .D(n2445), .CK(clk), .RN(n1553), .Q(
        \gbuff[11][21] ) );
  DFFRX1 \gbuff_reg[11][20]  ( .D(n2446), .CK(clk), .RN(n1553), .Q(
        \gbuff[11][20] ) );
  DFFRX1 \gbuff_reg[11][19]  ( .D(n2447), .CK(clk), .RN(n1552), .Q(
        \gbuff[11][19] ) );
  DFFRX1 \gbuff_reg[11][18]  ( .D(n2448), .CK(clk), .RN(n1552), .Q(
        \gbuff[11][18] ) );
  DFFRX1 \gbuff_reg[11][17]  ( .D(n2449), .CK(clk), .RN(n1552), .Q(
        \gbuff[11][17] ) );
  DFFRX1 \gbuff_reg[11][16]  ( .D(n2450), .CK(clk), .RN(n1552), .Q(
        \gbuff[11][16] ) );
  DFFRX1 \gbuff_reg[11][15]  ( .D(n2451), .CK(clk), .RN(n1552), .Q(
        \gbuff[11][15] ) );
  DFFRX1 \gbuff_reg[11][14]  ( .D(n2452), .CK(clk), .RN(n1552), .Q(
        \gbuff[11][14] ) );
  DFFRX1 \gbuff_reg[11][13]  ( .D(n2453), .CK(clk), .RN(n1552), .Q(
        \gbuff[11][13] ) );
  DFFRX1 \gbuff_reg[11][12]  ( .D(n2454), .CK(clk), .RN(n1552), .Q(
        \gbuff[11][12] ) );
  DFFRX1 \gbuff_reg[11][11]  ( .D(n2455), .CK(clk), .RN(n1552), .Q(
        \gbuff[11][11] ) );
  DFFRX1 \gbuff_reg[11][10]  ( .D(n2456), .CK(clk), .RN(n1552), .Q(
        \gbuff[11][10] ) );
  DFFRX1 \gbuff_reg[11][9]  ( .D(n2457), .CK(clk), .RN(n1552), .Q(
        \gbuff[11][9] ) );
  DFFRX1 \gbuff_reg[11][8]  ( .D(n2458), .CK(clk), .RN(n1552), .Q(
        \gbuff[11][8] ) );
  DFFRX1 \gbuff_reg[11][7]  ( .D(n2459), .CK(clk), .RN(n1551), .Q(
        \gbuff[11][7] ) );
  DFFRX1 \gbuff_reg[11][6]  ( .D(n2460), .CK(clk), .RN(n1551), .Q(
        \gbuff[11][6] ) );
  DFFRX1 \gbuff_reg[11][5]  ( .D(n2461), .CK(clk), .RN(n1551), .Q(
        \gbuff[11][5] ) );
  DFFRX1 \gbuff_reg[11][4]  ( .D(n2462), .CK(clk), .RN(n1551), .Q(
        \gbuff[11][4] ) );
  DFFRX1 \gbuff_reg[11][3]  ( .D(n2463), .CK(clk), .RN(n1551), .Q(
        \gbuff[11][3] ) );
  DFFRX1 \gbuff_reg[11][2]  ( .D(n2464), .CK(clk), .RN(n1551), .Q(
        \gbuff[11][2] ) );
  DFFRX1 \gbuff_reg[11][1]  ( .D(n2465), .CK(clk), .RN(n1551), .Q(
        \gbuff[11][1] ) );
  DFFRX1 \gbuff_reg[11][0]  ( .D(n2466), .CK(clk), .RN(n1551), .Q(
        \gbuff[11][0] ) );
  DFFRX1 \gbuff_reg[7][31]  ( .D(n2563), .CK(clk), .RN(n1543), .Q(
        \gbuff[7][31] ) );
  DFFRX1 \gbuff_reg[7][30]  ( .D(n2564), .CK(clk), .RN(n1543), .Q(
        \gbuff[7][30] ) );
  DFFRX1 \gbuff_reg[7][29]  ( .D(n2565), .CK(clk), .RN(n1543), .Q(
        \gbuff[7][29] ) );
  DFFRX1 \gbuff_reg[7][28]  ( .D(n2566), .CK(clk), .RN(n1543), .Q(
        \gbuff[7][28] ) );
  DFFRX1 \gbuff_reg[7][27]  ( .D(n2567), .CK(clk), .RN(n1542), .Q(
        \gbuff[7][27] ) );
  DFFRX1 \gbuff_reg[7][26]  ( .D(n2568), .CK(clk), .RN(n1542), .Q(
        \gbuff[7][26] ) );
  DFFRX1 \gbuff_reg[7][25]  ( .D(n2569), .CK(clk), .RN(n1542), .Q(
        \gbuff[7][25] ) );
  DFFRX1 \gbuff_reg[7][24]  ( .D(n2570), .CK(clk), .RN(n1542), .Q(
        \gbuff[7][24] ) );
  DFFRX1 \gbuff_reg[7][23]  ( .D(n2571), .CK(clk), .RN(n1542), .Q(
        \gbuff[7][23] ) );
  DFFRX1 \gbuff_reg[7][22]  ( .D(n2572), .CK(clk), .RN(n1542), .Q(
        \gbuff[7][22] ) );
  DFFRX1 \gbuff_reg[7][21]  ( .D(n2573), .CK(clk), .RN(n1542), .Q(
        \gbuff[7][21] ) );
  DFFRX1 \gbuff_reg[7][20]  ( .D(n2574), .CK(clk), .RN(n1542), .Q(
        \gbuff[7][20] ) );
  DFFRX1 \gbuff_reg[7][19]  ( .D(n2575), .CK(clk), .RN(n1542), .Q(
        \gbuff[7][19] ) );
  DFFRX1 \gbuff_reg[7][18]  ( .D(n2576), .CK(clk), .RN(n1542), .Q(
        \gbuff[7][18] ) );
  DFFRX1 \gbuff_reg[7][17]  ( .D(n2577), .CK(clk), .RN(n1542), .Q(
        \gbuff[7][17] ) );
  DFFRX1 \gbuff_reg[7][16]  ( .D(n2578), .CK(clk), .RN(n1542), .Q(
        \gbuff[7][16] ) );
  DFFRX1 \gbuff_reg[7][15]  ( .D(n2579), .CK(clk), .RN(n1541), .Q(
        \gbuff[7][15] ) );
  DFFRX1 \gbuff_reg[7][14]  ( .D(n2580), .CK(clk), .RN(n1541), .Q(
        \gbuff[7][14] ) );
  DFFRX1 \gbuff_reg[7][13]  ( .D(n2581), .CK(clk), .RN(n1541), .Q(
        \gbuff[7][13] ) );
  DFFRX1 \gbuff_reg[7][12]  ( .D(n2582), .CK(clk), .RN(n1541), .Q(
        \gbuff[7][12] ) );
  DFFRX1 \gbuff_reg[7][11]  ( .D(n2583), .CK(clk), .RN(n1541), .Q(
        \gbuff[7][11] ) );
  DFFRX1 \gbuff_reg[7][10]  ( .D(n2584), .CK(clk), .RN(n1541), .Q(
        \gbuff[7][10] ) );
  DFFRX1 \gbuff_reg[7][9]  ( .D(n2585), .CK(clk), .RN(n1541), .Q(\gbuff[7][9] ) );
  DFFRX1 \gbuff_reg[7][8]  ( .D(n2586), .CK(clk), .RN(n1541), .Q(\gbuff[7][8] ) );
  DFFRX1 \gbuff_reg[7][7]  ( .D(n2587), .CK(clk), .RN(n1541), .Q(\gbuff[7][7] ) );
  DFFRX1 \gbuff_reg[7][6]  ( .D(n2588), .CK(clk), .RN(n1541), .Q(\gbuff[7][6] ) );
  DFFRX1 \gbuff_reg[7][5]  ( .D(n2589), .CK(clk), .RN(n1541), .Q(\gbuff[7][5] ) );
  DFFRX1 \gbuff_reg[7][4]  ( .D(n2590), .CK(clk), .RN(n1541), .Q(\gbuff[7][4] ) );
  DFFRX1 \gbuff_reg[7][3]  ( .D(n2591), .CK(clk), .RN(n1540), .Q(\gbuff[7][3] ) );
  DFFRX1 \gbuff_reg[7][2]  ( .D(n2592), .CK(clk), .RN(n1540), .Q(\gbuff[7][2] ) );
  DFFRX1 \gbuff_reg[7][1]  ( .D(n2593), .CK(clk), .RN(n1540), .Q(\gbuff[7][1] ) );
  DFFRX1 \gbuff_reg[7][0]  ( .D(n2594), .CK(clk), .RN(n1540), .Q(\gbuff[7][0] ) );
  DFFRX1 \gbuff_reg[3][31]  ( .D(n2691), .CK(clk), .RN(n1532), .Q(
        \gbuff[3][31] ) );
  DFFRX1 \gbuff_reg[3][30]  ( .D(n2692), .CK(clk), .RN(n1532), .Q(
        \gbuff[3][30] ) );
  DFFRX1 \gbuff_reg[3][29]  ( .D(n2693), .CK(clk), .RN(n1532), .Q(
        \gbuff[3][29] ) );
  DFFRX1 \gbuff_reg[3][28]  ( .D(n2694), .CK(clk), .RN(n1532), .Q(
        \gbuff[3][28] ) );
  DFFRX1 \gbuff_reg[3][27]  ( .D(n2695), .CK(clk), .RN(n1532), .Q(
        \gbuff[3][27] ) );
  DFFRX1 \gbuff_reg[3][26]  ( .D(n2696), .CK(clk), .RN(n1532), .Q(
        \gbuff[3][26] ) );
  DFFRX1 \gbuff_reg[3][25]  ( .D(n2697), .CK(clk), .RN(n1532), .Q(
        \gbuff[3][25] ) );
  DFFRX1 \gbuff_reg[3][24]  ( .D(n2698), .CK(clk), .RN(n1532), .Q(
        \gbuff[3][24] ) );
  DFFRX1 \gbuff_reg[3][23]  ( .D(n2699), .CK(clk), .RN(n1531), .Q(
        \gbuff[3][23] ) );
  DFFRX1 \gbuff_reg[3][22]  ( .D(n2700), .CK(clk), .RN(n1531), .Q(
        \gbuff[3][22] ) );
  DFFRX1 \gbuff_reg[3][21]  ( .D(n2701), .CK(clk), .RN(n1531), .Q(
        \gbuff[3][21] ) );
  DFFRX1 \gbuff_reg[3][20]  ( .D(n2702), .CK(clk), .RN(n1531), .Q(
        \gbuff[3][20] ) );
  DFFRX1 \gbuff_reg[3][19]  ( .D(n2703), .CK(clk), .RN(n1531), .Q(
        \gbuff[3][19] ) );
  DFFRX1 \gbuff_reg[3][18]  ( .D(n2704), .CK(clk), .RN(n1531), .Q(
        \gbuff[3][18] ) );
  DFFRX1 \gbuff_reg[3][17]  ( .D(n2705), .CK(clk), .RN(n1531), .Q(
        \gbuff[3][17] ) );
  DFFRX1 \gbuff_reg[3][16]  ( .D(n2706), .CK(clk), .RN(n1531), .Q(
        \gbuff[3][16] ) );
  DFFRX1 \gbuff_reg[3][15]  ( .D(n2707), .CK(clk), .RN(n1531), .Q(
        \gbuff[3][15] ) );
  DFFRX1 \gbuff_reg[3][14]  ( .D(n2708), .CK(clk), .RN(n1531), .Q(
        \gbuff[3][14] ) );
  DFFRX1 \gbuff_reg[3][13]  ( .D(n2709), .CK(clk), .RN(n1531), .Q(
        \gbuff[3][13] ) );
  DFFRX1 \gbuff_reg[3][12]  ( .D(n2710), .CK(clk), .RN(n1531), .Q(
        \gbuff[3][12] ) );
  DFFRX1 \gbuff_reg[3][11]  ( .D(n2711), .CK(clk), .RN(n1530), .Q(
        \gbuff[3][11] ) );
  DFFRX1 \gbuff_reg[3][10]  ( .D(n2712), .CK(clk), .RN(n1530), .Q(
        \gbuff[3][10] ) );
  DFFRX1 \gbuff_reg[3][9]  ( .D(n2713), .CK(clk), .RN(n1530), .Q(\gbuff[3][9] ) );
  DFFRX1 \gbuff_reg[3][8]  ( .D(n2714), .CK(clk), .RN(n1530), .Q(\gbuff[3][8] ) );
  DFFRX1 \gbuff_reg[3][7]  ( .D(n2715), .CK(clk), .RN(n1530), .Q(\gbuff[3][7] ) );
  DFFRX1 \gbuff_reg[3][6]  ( .D(n2716), .CK(clk), .RN(n1530), .Q(\gbuff[3][6] ) );
  DFFRX1 \gbuff_reg[3][5]  ( .D(n2717), .CK(clk), .RN(n1530), .Q(\gbuff[3][5] ) );
  DFFRX1 \gbuff_reg[3][4]  ( .D(n2718), .CK(clk), .RN(n1530), .Q(\gbuff[3][4] ) );
  DFFRX1 \gbuff_reg[3][3]  ( .D(n2719), .CK(clk), .RN(n1530), .Q(\gbuff[3][3] ) );
  DFFRX1 \gbuff_reg[3][2]  ( .D(n2720), .CK(clk), .RN(n1530), .Q(\gbuff[3][2] ) );
  DFFRX1 \gbuff_reg[3][1]  ( .D(n2721), .CK(clk), .RN(n1530), .Q(\gbuff[3][1] ) );
  DFFRX1 \gbuff_reg[3][0]  ( .D(n2722), .CK(clk), .RN(n1530), .Q(\gbuff[3][0] ) );
  DFFRX1 \gbuff_reg[28][31]  ( .D(n1891), .CK(clk), .RN(n1599), .Q(
        \gbuff[28][31] ) );
  DFFRX1 \gbuff_reg[28][30]  ( .D(n1892), .CK(clk), .RN(n1599), .Q(
        \gbuff[28][30] ) );
  DFFRX1 \gbuff_reg[28][29]  ( .D(n1893), .CK(clk), .RN(n1599), .Q(
        \gbuff[28][29] ) );
  DFFRX1 \gbuff_reg[28][28]  ( .D(n1894), .CK(clk), .RN(n1599), .Q(
        \gbuff[28][28] ) );
  DFFRX1 \gbuff_reg[28][27]  ( .D(n1895), .CK(clk), .RN(n1598), .Q(
        \gbuff[28][27] ) );
  DFFRX1 \gbuff_reg[28][26]  ( .D(n1896), .CK(clk), .RN(n1598), .Q(
        \gbuff[28][26] ) );
  DFFRX1 \gbuff_reg[28][25]  ( .D(n1897), .CK(clk), .RN(n1598), .Q(
        \gbuff[28][25] ) );
  DFFRX1 \gbuff_reg[28][24]  ( .D(n1898), .CK(clk), .RN(n1598), .Q(
        \gbuff[28][24] ) );
  DFFRX1 \gbuff_reg[28][23]  ( .D(n1899), .CK(clk), .RN(n1598), .Q(
        \gbuff[28][23] ) );
  DFFRX1 \gbuff_reg[28][22]  ( .D(n1900), .CK(clk), .RN(n1598), .Q(
        \gbuff[28][22] ) );
  DFFRX1 \gbuff_reg[28][21]  ( .D(n1901), .CK(clk), .RN(n1598), .Q(
        \gbuff[28][21] ) );
  DFFRX1 \gbuff_reg[28][20]  ( .D(n1902), .CK(clk), .RN(n1598), .Q(
        \gbuff[28][20] ) );
  DFFRX1 \gbuff_reg[28][19]  ( .D(n1903), .CK(clk), .RN(n1598), .Q(
        \gbuff[28][19] ) );
  DFFRX1 \gbuff_reg[28][18]  ( .D(n1904), .CK(clk), .RN(n1598), .Q(
        \gbuff[28][18] ) );
  DFFRX1 \gbuff_reg[28][17]  ( .D(n1905), .CK(clk), .RN(n1598), .Q(
        \gbuff[28][17] ) );
  DFFRX1 \gbuff_reg[28][16]  ( .D(n1906), .CK(clk), .RN(n1598), .Q(
        \gbuff[28][16] ) );
  DFFRX1 \gbuff_reg[28][15]  ( .D(n1907), .CK(clk), .RN(n1597), .Q(
        \gbuff[28][15] ) );
  DFFRX1 \gbuff_reg[28][14]  ( .D(n1908), .CK(clk), .RN(n1597), .Q(
        \gbuff[28][14] ) );
  DFFRX1 \gbuff_reg[28][13]  ( .D(n1909), .CK(clk), .RN(n1597), .Q(
        \gbuff[28][13] ) );
  DFFRX1 \gbuff_reg[28][12]  ( .D(n1910), .CK(clk), .RN(n1597), .Q(
        \gbuff[28][12] ) );
  DFFRX1 \gbuff_reg[28][11]  ( .D(n1911), .CK(clk), .RN(n1597), .Q(
        \gbuff[28][11] ) );
  DFFRX1 \gbuff_reg[28][10]  ( .D(n1912), .CK(clk), .RN(n1597), .Q(
        \gbuff[28][10] ) );
  DFFRX1 \gbuff_reg[28][9]  ( .D(n1913), .CK(clk), .RN(n1597), .Q(
        \gbuff[28][9] ) );
  DFFRX1 \gbuff_reg[28][8]  ( .D(n1914), .CK(clk), .RN(n1597), .Q(
        \gbuff[28][8] ) );
  DFFRX1 \gbuff_reg[28][7]  ( .D(n1915), .CK(clk), .RN(n1597), .Q(
        \gbuff[28][7] ) );
  DFFRX1 \gbuff_reg[28][6]  ( .D(n1916), .CK(clk), .RN(n1597), .Q(
        \gbuff[28][6] ) );
  DFFRX1 \gbuff_reg[28][5]  ( .D(n1917), .CK(clk), .RN(n1597), .Q(
        \gbuff[28][5] ) );
  DFFRX1 \gbuff_reg[28][4]  ( .D(n1918), .CK(clk), .RN(n1597), .Q(
        \gbuff[28][4] ) );
  DFFRX1 \gbuff_reg[28][3]  ( .D(n1919), .CK(clk), .RN(n1596), .Q(
        \gbuff[28][3] ) );
  DFFRX1 \gbuff_reg[28][2]  ( .D(n1920), .CK(clk), .RN(n1596), .Q(
        \gbuff[28][2] ) );
  DFFRX1 \gbuff_reg[28][1]  ( .D(n1921), .CK(clk), .RN(n1596), .Q(
        \gbuff[28][1] ) );
  DFFRX1 \gbuff_reg[28][0]  ( .D(n1922), .CK(clk), .RN(n1596), .Q(
        \gbuff[28][0] ) );
  DFFRX1 \gbuff_reg[24][31]  ( .D(n2019), .CK(clk), .RN(n1588), .Q(
        \gbuff[24][31] ) );
  DFFRX1 \gbuff_reg[24][30]  ( .D(n2020), .CK(clk), .RN(n1588), .Q(
        \gbuff[24][30] ) );
  DFFRX1 \gbuff_reg[24][29]  ( .D(n2021), .CK(clk), .RN(n1588), .Q(
        \gbuff[24][29] ) );
  DFFRX1 \gbuff_reg[24][28]  ( .D(n2022), .CK(clk), .RN(n1588), .Q(
        \gbuff[24][28] ) );
  DFFRX1 \gbuff_reg[24][27]  ( .D(n2023), .CK(clk), .RN(n1588), .Q(
        \gbuff[24][27] ) );
  DFFRX1 \gbuff_reg[24][26]  ( .D(n2024), .CK(clk), .RN(n1588), .Q(
        \gbuff[24][26] ) );
  DFFRX1 \gbuff_reg[24][25]  ( .D(n2025), .CK(clk), .RN(n1588), .Q(
        \gbuff[24][25] ) );
  DFFRX1 \gbuff_reg[24][24]  ( .D(n2026), .CK(clk), .RN(n1588), .Q(
        \gbuff[24][24] ) );
  DFFRX1 \gbuff_reg[24][23]  ( .D(n2027), .CK(clk), .RN(n1587), .Q(
        \gbuff[24][23] ) );
  DFFRX1 \gbuff_reg[24][22]  ( .D(n2028), .CK(clk), .RN(n1587), .Q(
        \gbuff[24][22] ) );
  DFFRX1 \gbuff_reg[24][21]  ( .D(n2029), .CK(clk), .RN(n1587), .Q(
        \gbuff[24][21] ) );
  DFFRX1 \gbuff_reg[24][20]  ( .D(n2030), .CK(clk), .RN(n1587), .Q(
        \gbuff[24][20] ) );
  DFFRX1 \gbuff_reg[24][19]  ( .D(n2031), .CK(clk), .RN(n1587), .Q(
        \gbuff[24][19] ) );
  DFFRX1 \gbuff_reg[24][18]  ( .D(n2032), .CK(clk), .RN(n1587), .Q(
        \gbuff[24][18] ) );
  DFFRX1 \gbuff_reg[24][17]  ( .D(n2033), .CK(clk), .RN(n1587), .Q(
        \gbuff[24][17] ) );
  DFFRX1 \gbuff_reg[24][16]  ( .D(n2034), .CK(clk), .RN(n1587), .Q(
        \gbuff[24][16] ) );
  DFFRX1 \gbuff_reg[24][15]  ( .D(n2035), .CK(clk), .RN(n1587), .Q(
        \gbuff[24][15] ) );
  DFFRX1 \gbuff_reg[24][14]  ( .D(n2036), .CK(clk), .RN(n1587), .Q(
        \gbuff[24][14] ) );
  DFFRX1 \gbuff_reg[24][13]  ( .D(n2037), .CK(clk), .RN(n1587), .Q(
        \gbuff[24][13] ) );
  DFFRX1 \gbuff_reg[24][12]  ( .D(n2038), .CK(clk), .RN(n1587), .Q(
        \gbuff[24][12] ) );
  DFFRX1 \gbuff_reg[24][11]  ( .D(n2039), .CK(clk), .RN(n1586), .Q(
        \gbuff[24][11] ) );
  DFFRX1 \gbuff_reg[24][10]  ( .D(n2040), .CK(clk), .RN(n1586), .Q(
        \gbuff[24][10] ) );
  DFFRX1 \gbuff_reg[24][9]  ( .D(n2041), .CK(clk), .RN(n1586), .Q(
        \gbuff[24][9] ) );
  DFFRX1 \gbuff_reg[24][8]  ( .D(n2042), .CK(clk), .RN(n1586), .Q(
        \gbuff[24][8] ) );
  DFFRX1 \gbuff_reg[24][7]  ( .D(n2043), .CK(clk), .RN(n1586), .Q(
        \gbuff[24][7] ) );
  DFFRX1 \gbuff_reg[24][6]  ( .D(n2044), .CK(clk), .RN(n1586), .Q(
        \gbuff[24][6] ) );
  DFFRX1 \gbuff_reg[24][5]  ( .D(n2045), .CK(clk), .RN(n1586), .Q(
        \gbuff[24][5] ) );
  DFFRX1 \gbuff_reg[24][4]  ( .D(n2046), .CK(clk), .RN(n1586), .Q(
        \gbuff[24][4] ) );
  DFFRX1 \gbuff_reg[24][3]  ( .D(n2047), .CK(clk), .RN(n1586), .Q(
        \gbuff[24][3] ) );
  DFFRX1 \gbuff_reg[24][2]  ( .D(n2048), .CK(clk), .RN(n1586), .Q(
        \gbuff[24][2] ) );
  DFFRX1 \gbuff_reg[24][1]  ( .D(n2049), .CK(clk), .RN(n1586), .Q(
        \gbuff[24][1] ) );
  DFFRX1 \gbuff_reg[24][0]  ( .D(n2050), .CK(clk), .RN(n1586), .Q(
        \gbuff[24][0] ) );
  DFFRX1 \gbuff_reg[20][31]  ( .D(n2147), .CK(clk), .RN(n1577), .Q(
        \gbuff[20][31] ) );
  DFFRX1 \gbuff_reg[20][30]  ( .D(n2148), .CK(clk), .RN(n1577), .Q(
        \gbuff[20][30] ) );
  DFFRX1 \gbuff_reg[20][29]  ( .D(n2149), .CK(clk), .RN(n1577), .Q(
        \gbuff[20][29] ) );
  DFFRX1 \gbuff_reg[20][28]  ( .D(n2150), .CK(clk), .RN(n1577), .Q(
        \gbuff[20][28] ) );
  DFFRX1 \gbuff_reg[20][27]  ( .D(n2151), .CK(clk), .RN(n1577), .Q(
        \gbuff[20][27] ) );
  DFFRX1 \gbuff_reg[20][26]  ( .D(n2152), .CK(clk), .RN(n1577), .Q(
        \gbuff[20][26] ) );
  DFFRX1 \gbuff_reg[20][25]  ( .D(n2153), .CK(clk), .RN(n1577), .Q(
        \gbuff[20][25] ) );
  DFFRX1 \gbuff_reg[20][24]  ( .D(n2154), .CK(clk), .RN(n1577), .Q(
        \gbuff[20][24] ) );
  DFFRX1 \gbuff_reg[20][23]  ( .D(n2155), .CK(clk), .RN(n1577), .Q(
        \gbuff[20][23] ) );
  DFFRX1 \gbuff_reg[20][22]  ( .D(n2156), .CK(clk), .RN(n1577), .Q(
        \gbuff[20][22] ) );
  DFFRX1 \gbuff_reg[20][21]  ( .D(n2157), .CK(clk), .RN(n1577), .Q(
        \gbuff[20][21] ) );
  DFFRX1 \gbuff_reg[20][20]  ( .D(n2158), .CK(clk), .RN(n1577), .Q(
        \gbuff[20][20] ) );
  DFFRX1 \gbuff_reg[20][19]  ( .D(n2159), .CK(clk), .RN(n1576), .Q(
        \gbuff[20][19] ) );
  DFFRX1 \gbuff_reg[20][18]  ( .D(n2160), .CK(clk), .RN(n1576), .Q(
        \gbuff[20][18] ) );
  DFFRX1 \gbuff_reg[20][17]  ( .D(n2161), .CK(clk), .RN(n1576), .Q(
        \gbuff[20][17] ) );
  DFFRX1 \gbuff_reg[20][16]  ( .D(n2162), .CK(clk), .RN(n1576), .Q(
        \gbuff[20][16] ) );
  DFFRX1 \gbuff_reg[20][15]  ( .D(n2163), .CK(clk), .RN(n1576), .Q(
        \gbuff[20][15] ) );
  DFFRX1 \gbuff_reg[20][14]  ( .D(n2164), .CK(clk), .RN(n1576), .Q(
        \gbuff[20][14] ) );
  DFFRX1 \gbuff_reg[20][13]  ( .D(n2165), .CK(clk), .RN(n1576), .Q(
        \gbuff[20][13] ) );
  DFFRX1 \gbuff_reg[20][12]  ( .D(n2166), .CK(clk), .RN(n1576), .Q(
        \gbuff[20][12] ) );
  DFFRX1 \gbuff_reg[20][11]  ( .D(n2167), .CK(clk), .RN(n1576), .Q(
        \gbuff[20][11] ) );
  DFFRX1 \gbuff_reg[20][10]  ( .D(n2168), .CK(clk), .RN(n1576), .Q(
        \gbuff[20][10] ) );
  DFFRX1 \gbuff_reg[20][9]  ( .D(n2169), .CK(clk), .RN(n1576), .Q(
        \gbuff[20][9] ) );
  DFFRX1 \gbuff_reg[20][8]  ( .D(n2170), .CK(clk), .RN(n1576), .Q(
        \gbuff[20][8] ) );
  DFFRX1 \gbuff_reg[20][7]  ( .D(n2171), .CK(clk), .RN(n1575), .Q(
        \gbuff[20][7] ) );
  DFFRX1 \gbuff_reg[20][6]  ( .D(n2172), .CK(clk), .RN(n1575), .Q(
        \gbuff[20][6] ) );
  DFFRX1 \gbuff_reg[20][5]  ( .D(n2173), .CK(clk), .RN(n1575), .Q(
        \gbuff[20][5] ) );
  DFFRX1 \gbuff_reg[20][4]  ( .D(n2174), .CK(clk), .RN(n1575), .Q(
        \gbuff[20][4] ) );
  DFFRX1 \gbuff_reg[20][3]  ( .D(n2175), .CK(clk), .RN(n1575), .Q(
        \gbuff[20][3] ) );
  DFFRX1 \gbuff_reg[20][2]  ( .D(n2176), .CK(clk), .RN(n1575), .Q(
        \gbuff[20][2] ) );
  DFFRX1 \gbuff_reg[20][1]  ( .D(n2177), .CK(clk), .RN(n1575), .Q(
        \gbuff[20][1] ) );
  DFFRX1 \gbuff_reg[20][0]  ( .D(n2178), .CK(clk), .RN(n1575), .Q(
        \gbuff[20][0] ) );
  DFFRX1 \gbuff_reg[16][31]  ( .D(n2275), .CK(clk), .RN(n1567), .Q(
        \gbuff[16][31] ) );
  DFFRX1 \gbuff_reg[16][30]  ( .D(n2276), .CK(clk), .RN(n1567), .Q(
        \gbuff[16][30] ) );
  DFFRX1 \gbuff_reg[16][29]  ( .D(n2277), .CK(clk), .RN(n1567), .Q(
        \gbuff[16][29] ) );
  DFFRX1 \gbuff_reg[16][28]  ( .D(n2278), .CK(clk), .RN(n1567), .Q(
        \gbuff[16][28] ) );
  DFFRX1 \gbuff_reg[16][27]  ( .D(n2279), .CK(clk), .RN(n1566), .Q(
        \gbuff[16][27] ) );
  DFFRX1 \gbuff_reg[16][26]  ( .D(n2280), .CK(clk), .RN(n1566), .Q(
        \gbuff[16][26] ) );
  DFFRX1 \gbuff_reg[16][25]  ( .D(n2281), .CK(clk), .RN(n1566), .Q(
        \gbuff[16][25] ) );
  DFFRX1 \gbuff_reg[16][24]  ( .D(n2282), .CK(clk), .RN(n1566), .Q(
        \gbuff[16][24] ) );
  DFFRX1 \gbuff_reg[16][23]  ( .D(n2283), .CK(clk), .RN(n1566), .Q(
        \gbuff[16][23] ) );
  DFFRX1 \gbuff_reg[16][22]  ( .D(n2284), .CK(clk), .RN(n1566), .Q(
        \gbuff[16][22] ) );
  DFFRX1 \gbuff_reg[16][21]  ( .D(n2285), .CK(clk), .RN(n1566), .Q(
        \gbuff[16][21] ) );
  DFFRX1 \gbuff_reg[16][20]  ( .D(n2286), .CK(clk), .RN(n1566), .Q(
        \gbuff[16][20] ) );
  DFFRX1 \gbuff_reg[16][19]  ( .D(n2287), .CK(clk), .RN(n1566), .Q(
        \gbuff[16][19] ) );
  DFFRX1 \gbuff_reg[16][18]  ( .D(n2288), .CK(clk), .RN(n1566), .Q(
        \gbuff[16][18] ) );
  DFFRX1 \gbuff_reg[16][17]  ( .D(n2289), .CK(clk), .RN(n1566), .Q(
        \gbuff[16][17] ) );
  DFFRX1 \gbuff_reg[16][16]  ( .D(n2290), .CK(clk), .RN(n1566), .Q(
        \gbuff[16][16] ) );
  DFFRX1 \gbuff_reg[16][15]  ( .D(n2291), .CK(clk), .RN(n1565), .Q(
        \gbuff[16][15] ) );
  DFFRX1 \gbuff_reg[16][14]  ( .D(n2292), .CK(clk), .RN(n1565), .Q(
        \gbuff[16][14] ) );
  DFFRX1 \gbuff_reg[16][13]  ( .D(n2293), .CK(clk), .RN(n1565), .Q(
        \gbuff[16][13] ) );
  DFFRX1 \gbuff_reg[16][12]  ( .D(n2294), .CK(clk), .RN(n1565), .Q(
        \gbuff[16][12] ) );
  DFFRX1 \gbuff_reg[16][11]  ( .D(n2295), .CK(clk), .RN(n1565), .Q(
        \gbuff[16][11] ) );
  DFFRX1 \gbuff_reg[16][10]  ( .D(n2296), .CK(clk), .RN(n1565), .Q(
        \gbuff[16][10] ) );
  DFFRX1 \gbuff_reg[16][9]  ( .D(n2297), .CK(clk), .RN(n1565), .Q(
        \gbuff[16][9] ) );
  DFFRX1 \gbuff_reg[16][8]  ( .D(n2298), .CK(clk), .RN(n1565), .Q(
        \gbuff[16][8] ) );
  DFFRX1 \gbuff_reg[16][7]  ( .D(n2299), .CK(clk), .RN(n1565), .Q(
        \gbuff[16][7] ) );
  DFFRX1 \gbuff_reg[16][6]  ( .D(n2300), .CK(clk), .RN(n1565), .Q(
        \gbuff[16][6] ) );
  DFFRX1 \gbuff_reg[16][5]  ( .D(n2301), .CK(clk), .RN(n1565), .Q(
        \gbuff[16][5] ) );
  DFFRX1 \gbuff_reg[16][4]  ( .D(n2302), .CK(clk), .RN(n1565), .Q(
        \gbuff[16][4] ) );
  DFFRX1 \gbuff_reg[16][3]  ( .D(n2303), .CK(clk), .RN(n1564), .Q(
        \gbuff[16][3] ) );
  DFFRX1 \gbuff_reg[16][2]  ( .D(n2304), .CK(clk), .RN(n1564), .Q(
        \gbuff[16][2] ) );
  DFFRX1 \gbuff_reg[16][1]  ( .D(n2305), .CK(clk), .RN(n1564), .Q(
        \gbuff[16][1] ) );
  DFFRX1 \gbuff_reg[16][0]  ( .D(n2306), .CK(clk), .RN(n1564), .Q(
        \gbuff[16][0] ) );
  DFFRX1 \gbuff_reg[12][31]  ( .D(n2403), .CK(clk), .RN(n1556), .Q(
        \gbuff[12][31] ) );
  DFFRX1 \gbuff_reg[12][30]  ( .D(n2404), .CK(clk), .RN(n1556), .Q(
        \gbuff[12][30] ) );
  DFFRX1 \gbuff_reg[12][29]  ( .D(n2405), .CK(clk), .RN(n1556), .Q(
        \gbuff[12][29] ) );
  DFFRX1 \gbuff_reg[12][28]  ( .D(n2406), .CK(clk), .RN(n1556), .Q(
        \gbuff[12][28] ) );
  DFFRX1 \gbuff_reg[12][27]  ( .D(n2407), .CK(clk), .RN(n1556), .Q(
        \gbuff[12][27] ) );
  DFFRX1 \gbuff_reg[12][26]  ( .D(n2408), .CK(clk), .RN(n1556), .Q(
        \gbuff[12][26] ) );
  DFFRX1 \gbuff_reg[12][25]  ( .D(n2409), .CK(clk), .RN(n1556), .Q(
        \gbuff[12][25] ) );
  DFFRX1 \gbuff_reg[12][24]  ( .D(n2410), .CK(clk), .RN(n1556), .Q(
        \gbuff[12][24] ) );
  DFFRX1 \gbuff_reg[12][23]  ( .D(n2411), .CK(clk), .RN(n1555), .Q(
        \gbuff[12][23] ) );
  DFFRX1 \gbuff_reg[12][22]  ( .D(n2412), .CK(clk), .RN(n1555), .Q(
        \gbuff[12][22] ) );
  DFFRX1 \gbuff_reg[12][21]  ( .D(n2413), .CK(clk), .RN(n1555), .Q(
        \gbuff[12][21] ) );
  DFFRX1 \gbuff_reg[12][20]  ( .D(n2414), .CK(clk), .RN(n1555), .Q(
        \gbuff[12][20] ) );
  DFFRX1 \gbuff_reg[12][19]  ( .D(n2415), .CK(clk), .RN(n1555), .Q(
        \gbuff[12][19] ) );
  DFFRX1 \gbuff_reg[12][18]  ( .D(n2416), .CK(clk), .RN(n1555), .Q(
        \gbuff[12][18] ) );
  DFFRX1 \gbuff_reg[12][17]  ( .D(n2417), .CK(clk), .RN(n1555), .Q(
        \gbuff[12][17] ) );
  DFFRX1 \gbuff_reg[12][16]  ( .D(n2418), .CK(clk), .RN(n1555), .Q(
        \gbuff[12][16] ) );
  DFFRX1 \gbuff_reg[12][15]  ( .D(n2419), .CK(clk), .RN(n1555), .Q(
        \gbuff[12][15] ) );
  DFFRX1 \gbuff_reg[12][14]  ( .D(n2420), .CK(clk), .RN(n1555), .Q(
        \gbuff[12][14] ) );
  DFFRX1 \gbuff_reg[12][13]  ( .D(n2421), .CK(clk), .RN(n1555), .Q(
        \gbuff[12][13] ) );
  DFFRX1 \gbuff_reg[12][12]  ( .D(n2422), .CK(clk), .RN(n1555), .Q(
        \gbuff[12][12] ) );
  DFFRX1 \gbuff_reg[12][11]  ( .D(n2423), .CK(clk), .RN(n1554), .Q(
        \gbuff[12][11] ) );
  DFFRX1 \gbuff_reg[12][10]  ( .D(n2424), .CK(clk), .RN(n1554), .Q(
        \gbuff[12][10] ) );
  DFFRX1 \gbuff_reg[12][9]  ( .D(n2425), .CK(clk), .RN(n1554), .Q(
        \gbuff[12][9] ) );
  DFFRX1 \gbuff_reg[12][8]  ( .D(n2426), .CK(clk), .RN(n1554), .Q(
        \gbuff[12][8] ) );
  DFFRX1 \gbuff_reg[12][7]  ( .D(n2427), .CK(clk), .RN(n1554), .Q(
        \gbuff[12][7] ) );
  DFFRX1 \gbuff_reg[12][6]  ( .D(n2428), .CK(clk), .RN(n1554), .Q(
        \gbuff[12][6] ) );
  DFFRX1 \gbuff_reg[12][5]  ( .D(n2429), .CK(clk), .RN(n1554), .Q(
        \gbuff[12][5] ) );
  DFFRX1 \gbuff_reg[12][4]  ( .D(n2430), .CK(clk), .RN(n1554), .Q(
        \gbuff[12][4] ) );
  DFFRX1 \gbuff_reg[12][3]  ( .D(n2431), .CK(clk), .RN(n1554), .Q(
        \gbuff[12][3] ) );
  DFFRX1 \gbuff_reg[12][2]  ( .D(n2432), .CK(clk), .RN(n1554), .Q(
        \gbuff[12][2] ) );
  DFFRX1 \gbuff_reg[12][1]  ( .D(n2433), .CK(clk), .RN(n1554), .Q(
        \gbuff[12][1] ) );
  DFFRX1 \gbuff_reg[12][0]  ( .D(n2434), .CK(clk), .RN(n1554), .Q(
        \gbuff[12][0] ) );
  DFFRX1 \gbuff_reg[8][31]  ( .D(n2531), .CK(clk), .RN(n1545), .Q(
        \gbuff[8][31] ) );
  DFFRX1 \gbuff_reg[8][30]  ( .D(n2532), .CK(clk), .RN(n1545), .Q(
        \gbuff[8][30] ) );
  DFFRX1 \gbuff_reg[8][29]  ( .D(n2533), .CK(clk), .RN(n1545), .Q(
        \gbuff[8][29] ) );
  DFFRX1 \gbuff_reg[8][28]  ( .D(n2534), .CK(clk), .RN(n1545), .Q(
        \gbuff[8][28] ) );
  DFFRX1 \gbuff_reg[8][27]  ( .D(n2535), .CK(clk), .RN(n1545), .Q(
        \gbuff[8][27] ) );
  DFFRX1 \gbuff_reg[8][26]  ( .D(n2536), .CK(clk), .RN(n1545), .Q(
        \gbuff[8][26] ) );
  DFFRX1 \gbuff_reg[8][25]  ( .D(n2537), .CK(clk), .RN(n1545), .Q(
        \gbuff[8][25] ) );
  DFFRX1 \gbuff_reg[8][24]  ( .D(n2538), .CK(clk), .RN(n1545), .Q(
        \gbuff[8][24] ) );
  DFFRX1 \gbuff_reg[8][23]  ( .D(n2539), .CK(clk), .RN(n1545), .Q(
        \gbuff[8][23] ) );
  DFFRX1 \gbuff_reg[8][22]  ( .D(n2540), .CK(clk), .RN(n1545), .Q(
        \gbuff[8][22] ) );
  DFFRX1 \gbuff_reg[8][21]  ( .D(n2541), .CK(clk), .RN(n1545), .Q(
        \gbuff[8][21] ) );
  DFFRX1 \gbuff_reg[8][20]  ( .D(n2542), .CK(clk), .RN(n1545), .Q(
        \gbuff[8][20] ) );
  DFFRX1 \gbuff_reg[8][19]  ( .D(n2543), .CK(clk), .RN(n1544), .Q(
        \gbuff[8][19] ) );
  DFFRX1 \gbuff_reg[8][18]  ( .D(n2544), .CK(clk), .RN(n1544), .Q(
        \gbuff[8][18] ) );
  DFFRX1 \gbuff_reg[8][17]  ( .D(n2545), .CK(clk), .RN(n1544), .Q(
        \gbuff[8][17] ) );
  DFFRX1 \gbuff_reg[8][16]  ( .D(n2546), .CK(clk), .RN(n1544), .Q(
        \gbuff[8][16] ) );
  DFFRX1 \gbuff_reg[8][15]  ( .D(n2547), .CK(clk), .RN(n1544), .Q(
        \gbuff[8][15] ) );
  DFFRX1 \gbuff_reg[8][14]  ( .D(n2548), .CK(clk), .RN(n1544), .Q(
        \gbuff[8][14] ) );
  DFFRX1 \gbuff_reg[8][13]  ( .D(n2549), .CK(clk), .RN(n1544), .Q(
        \gbuff[8][13] ) );
  DFFRX1 \gbuff_reg[8][12]  ( .D(n2550), .CK(clk), .RN(n1544), .Q(
        \gbuff[8][12] ) );
  DFFRX1 \gbuff_reg[8][11]  ( .D(n2551), .CK(clk), .RN(n1544), .Q(
        \gbuff[8][11] ) );
  DFFRX1 \gbuff_reg[8][10]  ( .D(n2552), .CK(clk), .RN(n1544), .Q(
        \gbuff[8][10] ) );
  DFFRX1 \gbuff_reg[8][9]  ( .D(n2553), .CK(clk), .RN(n1544), .Q(\gbuff[8][9] ) );
  DFFRX1 \gbuff_reg[8][8]  ( .D(n2554), .CK(clk), .RN(n1544), .Q(\gbuff[8][8] ) );
  DFFRX1 \gbuff_reg[8][7]  ( .D(n2555), .CK(clk), .RN(n1543), .Q(\gbuff[8][7] ) );
  DFFRX1 \gbuff_reg[8][6]  ( .D(n2556), .CK(clk), .RN(n1543), .Q(\gbuff[8][6] ) );
  DFFRX1 \gbuff_reg[8][5]  ( .D(n2557), .CK(clk), .RN(n1543), .Q(\gbuff[8][5] ) );
  DFFRX1 \gbuff_reg[8][4]  ( .D(n2558), .CK(clk), .RN(n1543), .Q(\gbuff[8][4] ) );
  DFFRX1 \gbuff_reg[8][3]  ( .D(n2559), .CK(clk), .RN(n1543), .Q(\gbuff[8][3] ) );
  DFFRX1 \gbuff_reg[8][2]  ( .D(n2560), .CK(clk), .RN(n1543), .Q(\gbuff[8][2] ) );
  DFFRX1 \gbuff_reg[8][1]  ( .D(n2561), .CK(clk), .RN(n1543), .Q(\gbuff[8][1] ) );
  DFFRX1 \gbuff_reg[8][0]  ( .D(n2562), .CK(clk), .RN(n1543), .Q(\gbuff[8][0] ) );
  DFFRX1 \gbuff_reg[4][31]  ( .D(n2659), .CK(clk), .RN(n1535), .Q(
        \gbuff[4][31] ) );
  DFFRX1 \gbuff_reg[4][30]  ( .D(n2660), .CK(clk), .RN(n1535), .Q(
        \gbuff[4][30] ) );
  DFFRX1 \gbuff_reg[4][29]  ( .D(n2661), .CK(clk), .RN(n1535), .Q(
        \gbuff[4][29] ) );
  DFFRX1 \gbuff_reg[4][28]  ( .D(n2662), .CK(clk), .RN(n1535), .Q(
        \gbuff[4][28] ) );
  DFFRX1 \gbuff_reg[4][27]  ( .D(n2663), .CK(clk), .RN(n1534), .Q(
        \gbuff[4][27] ) );
  DFFRX1 \gbuff_reg[4][26]  ( .D(n2664), .CK(clk), .RN(n1534), .Q(
        \gbuff[4][26] ) );
  DFFRX1 \gbuff_reg[4][25]  ( .D(n2665), .CK(clk), .RN(n1534), .Q(
        \gbuff[4][25] ) );
  DFFRX1 \gbuff_reg[4][24]  ( .D(n2666), .CK(clk), .RN(n1534), .Q(
        \gbuff[4][24] ) );
  DFFRX1 \gbuff_reg[4][23]  ( .D(n2667), .CK(clk), .RN(n1534), .Q(
        \gbuff[4][23] ) );
  DFFRX1 \gbuff_reg[4][22]  ( .D(n2668), .CK(clk), .RN(n1534), .Q(
        \gbuff[4][22] ) );
  DFFRX1 \gbuff_reg[4][21]  ( .D(n2669), .CK(clk), .RN(n1534), .Q(
        \gbuff[4][21] ) );
  DFFRX1 \gbuff_reg[4][20]  ( .D(n2670), .CK(clk), .RN(n1534), .Q(
        \gbuff[4][20] ) );
  DFFRX1 \gbuff_reg[4][19]  ( .D(n2671), .CK(clk), .RN(n1534), .Q(
        \gbuff[4][19] ) );
  DFFRX1 \gbuff_reg[4][18]  ( .D(n2672), .CK(clk), .RN(n1534), .Q(
        \gbuff[4][18] ) );
  DFFRX1 \gbuff_reg[4][17]  ( .D(n2673), .CK(clk), .RN(n1534), .Q(
        \gbuff[4][17] ) );
  DFFRX1 \gbuff_reg[4][16]  ( .D(n2674), .CK(clk), .RN(n1534), .Q(
        \gbuff[4][16] ) );
  DFFRX1 \gbuff_reg[4][15]  ( .D(n2675), .CK(clk), .RN(n1533), .Q(
        \gbuff[4][15] ) );
  DFFRX1 \gbuff_reg[4][14]  ( .D(n2676), .CK(clk), .RN(n1533), .Q(
        \gbuff[4][14] ) );
  DFFRX1 \gbuff_reg[4][13]  ( .D(n2677), .CK(clk), .RN(n1533), .Q(
        \gbuff[4][13] ) );
  DFFRX1 \gbuff_reg[4][12]  ( .D(n2678), .CK(clk), .RN(n1533), .Q(
        \gbuff[4][12] ) );
  DFFRX1 \gbuff_reg[4][11]  ( .D(n2679), .CK(clk), .RN(n1533), .Q(
        \gbuff[4][11] ) );
  DFFRX1 \gbuff_reg[4][10]  ( .D(n2680), .CK(clk), .RN(n1533), .Q(
        \gbuff[4][10] ) );
  DFFRX1 \gbuff_reg[4][9]  ( .D(n2681), .CK(clk), .RN(n1533), .Q(\gbuff[4][9] ) );
  DFFRX1 \gbuff_reg[4][8]  ( .D(n2682), .CK(clk), .RN(n1533), .Q(\gbuff[4][8] ) );
  DFFRX1 \gbuff_reg[4][7]  ( .D(n2683), .CK(clk), .RN(n1533), .Q(\gbuff[4][7] ) );
  DFFRX1 \gbuff_reg[4][6]  ( .D(n2684), .CK(clk), .RN(n1533), .Q(\gbuff[4][6] ) );
  DFFRX1 \gbuff_reg[4][5]  ( .D(n2685), .CK(clk), .RN(n1533), .Q(\gbuff[4][5] ) );
  DFFRX1 \gbuff_reg[4][4]  ( .D(n2686), .CK(clk), .RN(n1533), .Q(\gbuff[4][4] ) );
  DFFRX1 \gbuff_reg[4][3]  ( .D(n2687), .CK(clk), .RN(n1532), .Q(\gbuff[4][3] ) );
  DFFRX1 \gbuff_reg[4][2]  ( .D(n2688), .CK(clk), .RN(n1532), .Q(\gbuff[4][2] ) );
  DFFRX1 \gbuff_reg[4][1]  ( .D(n2689), .CK(clk), .RN(n1532), .Q(\gbuff[4][1] ) );
  DFFRX1 \gbuff_reg[4][0]  ( .D(n2690), .CK(clk), .RN(n1532), .Q(\gbuff[4][0] ) );
  DFFRX1 \gbuff_reg[0][31]  ( .D(n2787), .CK(clk), .RN(n1524), .Q(
        \gbuff[0][31] ) );
  DFFRX1 \gbuff_reg[0][30]  ( .D(n2788), .CK(clk), .RN(n1524), .Q(
        \gbuff[0][30] ) );
  DFFRX1 \gbuff_reg[0][29]  ( .D(n2789), .CK(clk), .RN(n1524), .Q(
        \gbuff[0][29] ) );
  DFFRX1 \gbuff_reg[0][28]  ( .D(n2790), .CK(clk), .RN(n1524), .Q(
        \gbuff[0][28] ) );
  DFFRX1 \gbuff_reg[0][27]  ( .D(n2791), .CK(clk), .RN(n1524), .Q(
        \gbuff[0][27] ) );
  DFFRX1 \gbuff_reg[0][26]  ( .D(n2792), .CK(clk), .RN(n1524), .Q(
        \gbuff[0][26] ) );
  DFFRX1 \gbuff_reg[0][25]  ( .D(n2793), .CK(clk), .RN(n1524), .Q(
        \gbuff[0][25] ) );
  DFFRX1 \gbuff_reg[0][24]  ( .D(n2794), .CK(clk), .RN(n1524), .Q(
        \gbuff[0][24] ) );
  DFFRX1 \gbuff_reg[0][23]  ( .D(n2795), .CK(clk), .RN(n1523), .Q(
        \gbuff[0][23] ) );
  DFFRX1 \gbuff_reg[0][22]  ( .D(n2796), .CK(clk), .RN(n1523), .Q(
        \gbuff[0][22] ) );
  DFFRX1 \gbuff_reg[0][21]  ( .D(n2797), .CK(clk), .RN(n1523), .Q(
        \gbuff[0][21] ) );
  DFFRX1 \gbuff_reg[0][20]  ( .D(n2798), .CK(clk), .RN(n1523), .Q(
        \gbuff[0][20] ) );
  DFFRX1 \gbuff_reg[0][19]  ( .D(n2799), .CK(clk), .RN(n1523), .Q(
        \gbuff[0][19] ) );
  DFFRX1 \gbuff_reg[0][18]  ( .D(n2800), .CK(clk), .RN(n1523), .Q(
        \gbuff[0][18] ) );
  DFFRX1 \gbuff_reg[0][17]  ( .D(n2801), .CK(clk), .RN(n1523), .Q(
        \gbuff[0][17] ) );
  DFFRX1 \gbuff_reg[0][16]  ( .D(n2802), .CK(clk), .RN(n1523), .Q(
        \gbuff[0][16] ) );
  DFFRX1 \gbuff_reg[0][15]  ( .D(n2803), .CK(clk), .RN(n1523), .Q(
        \gbuff[0][15] ) );
  DFFRX1 \gbuff_reg[0][14]  ( .D(n2804), .CK(clk), .RN(n1523), .Q(
        \gbuff[0][14] ) );
  DFFRX1 \gbuff_reg[0][13]  ( .D(n2805), .CK(clk), .RN(n1523), .Q(
        \gbuff[0][13] ) );
  DFFRX1 \gbuff_reg[0][12]  ( .D(n2806), .CK(clk), .RN(n1523), .Q(
        \gbuff[0][12] ) );
  DFFRX1 \gbuff_reg[0][11]  ( .D(n2807), .CK(clk), .RN(n1522), .Q(
        \gbuff[0][11] ) );
  DFFRX1 \gbuff_reg[0][10]  ( .D(n2808), .CK(clk), .RN(n1522), .Q(
        \gbuff[0][10] ) );
  DFFRX1 \gbuff_reg[0][9]  ( .D(n2809), .CK(clk), .RN(n1522), .Q(\gbuff[0][9] ) );
  DFFRX1 \gbuff_reg[0][8]  ( .D(n2810), .CK(clk), .RN(n1522), .Q(\gbuff[0][8] ) );
  DFFRX1 \gbuff_reg[0][7]  ( .D(n2811), .CK(clk), .RN(n1522), .Q(\gbuff[0][7] ) );
  DFFRX1 \gbuff_reg[0][6]  ( .D(n2812), .CK(clk), .RN(n1522), .Q(\gbuff[0][6] ) );
  DFFRX1 \gbuff_reg[0][5]  ( .D(n2813), .CK(clk), .RN(n1522), .Q(\gbuff[0][5] ) );
  DFFRX1 \gbuff_reg[0][4]  ( .D(n2814), .CK(clk), .RN(n1522), .Q(\gbuff[0][4] ) );
  DFFRX1 \gbuff_reg[0][3]  ( .D(n2815), .CK(clk), .RN(n1522), .Q(\gbuff[0][3] ) );
  DFFRX1 \gbuff_reg[0][2]  ( .D(n2816), .CK(clk), .RN(n1522), .Q(\gbuff[0][2] ) );
  DFFRX1 \gbuff_reg[0][1]  ( .D(n2817), .CK(clk), .RN(n1522), .Q(\gbuff[0][1] ) );
  DFFRX1 \gbuff_reg[0][0]  ( .D(n2818), .CK(clk), .RN(n1522), .Q(\gbuff[0][0] ) );
  DFFRX1 \gbuff_reg[30][31]  ( .D(n1827), .CK(clk), .RN(n1604), .Q(
        \gbuff[30][31] ) );
  DFFRX1 \gbuff_reg[30][30]  ( .D(n1828), .CK(clk), .RN(n1604), .Q(
        \gbuff[30][30] ) );
  DFFRX1 \gbuff_reg[30][29]  ( .D(n1829), .CK(clk), .RN(n1604), .Q(
        \gbuff[30][29] ) );
  DFFRX1 \gbuff_reg[30][28]  ( .D(n1830), .CK(clk), .RN(n1604), .Q(
        \gbuff[30][28] ) );
  DFFRX1 \gbuff_reg[30][27]  ( .D(n1831), .CK(clk), .RN(n1604), .Q(
        \gbuff[30][27] ) );
  DFFRX1 \gbuff_reg[30][26]  ( .D(n1832), .CK(clk), .RN(n1604), .Q(
        \gbuff[30][26] ) );
  DFFRX1 \gbuff_reg[30][25]  ( .D(n1833), .CK(clk), .RN(n1604), .Q(
        \gbuff[30][25] ) );
  DFFRX1 \gbuff_reg[30][24]  ( .D(n1834), .CK(clk), .RN(n1604), .Q(
        \gbuff[30][24] ) );
  DFFRX1 \gbuff_reg[30][23]  ( .D(n1835), .CK(clk), .RN(n1603), .Q(
        \gbuff[30][23] ) );
  DFFRX1 \gbuff_reg[30][22]  ( .D(n1836), .CK(clk), .RN(n1603), .Q(
        \gbuff[30][22] ) );
  DFFRX1 \gbuff_reg[30][21]  ( .D(n1837), .CK(clk), .RN(n1603), .Q(
        \gbuff[30][21] ) );
  DFFRX1 \gbuff_reg[30][20]  ( .D(n1838), .CK(clk), .RN(n1603), .Q(
        \gbuff[30][20] ) );
  DFFRX1 \gbuff_reg[30][19]  ( .D(n1839), .CK(clk), .RN(n1603), .Q(
        \gbuff[30][19] ) );
  DFFRX1 \gbuff_reg[30][18]  ( .D(n1840), .CK(clk), .RN(n1603), .Q(
        \gbuff[30][18] ) );
  DFFRX1 \gbuff_reg[30][17]  ( .D(n1841), .CK(clk), .RN(n1603), .Q(
        \gbuff[30][17] ) );
  DFFRX1 \gbuff_reg[30][16]  ( .D(n1842), .CK(clk), .RN(n1603), .Q(
        \gbuff[30][16] ) );
  DFFRX1 \gbuff_reg[30][15]  ( .D(n1843), .CK(clk), .RN(n1603), .Q(
        \gbuff[30][15] ) );
  DFFRX1 \gbuff_reg[30][14]  ( .D(n1844), .CK(clk), .RN(n1603), .Q(
        \gbuff[30][14] ) );
  DFFRX1 \gbuff_reg[30][13]  ( .D(n1845), .CK(clk), .RN(n1603), .Q(
        \gbuff[30][13] ) );
  DFFRX1 \gbuff_reg[30][12]  ( .D(n1846), .CK(clk), .RN(n1603), .Q(
        \gbuff[30][12] ) );
  DFFRX1 \gbuff_reg[30][11]  ( .D(n1847), .CK(clk), .RN(n1602), .Q(
        \gbuff[30][11] ) );
  DFFRX1 \gbuff_reg[30][10]  ( .D(n1848), .CK(clk), .RN(n1602), .Q(
        \gbuff[30][10] ) );
  DFFRX1 \gbuff_reg[30][9]  ( .D(n1849), .CK(clk), .RN(n1602), .Q(
        \gbuff[30][9] ) );
  DFFRX1 \gbuff_reg[30][8]  ( .D(n1850), .CK(clk), .RN(n1602), .Q(
        \gbuff[30][8] ) );
  DFFRX1 \gbuff_reg[30][7]  ( .D(n1851), .CK(clk), .RN(n1602), .Q(
        \gbuff[30][7] ) );
  DFFRX1 \gbuff_reg[30][6]  ( .D(n1852), .CK(clk), .RN(n1602), .Q(
        \gbuff[30][6] ) );
  DFFRX1 \gbuff_reg[30][5]  ( .D(n1853), .CK(clk), .RN(n1602), .Q(
        \gbuff[30][5] ) );
  DFFRX1 \gbuff_reg[30][4]  ( .D(n1854), .CK(clk), .RN(n1602), .Q(
        \gbuff[30][4] ) );
  DFFRX1 \gbuff_reg[30][3]  ( .D(n1855), .CK(clk), .RN(n1602), .Q(
        \gbuff[30][3] ) );
  DFFRX1 \gbuff_reg[30][2]  ( .D(n1856), .CK(clk), .RN(n1602), .Q(
        \gbuff[30][2] ) );
  DFFRX1 \gbuff_reg[30][1]  ( .D(n1857), .CK(clk), .RN(n1602), .Q(
        \gbuff[30][1] ) );
  DFFRX1 \gbuff_reg[30][0]  ( .D(n1858), .CK(clk), .RN(n1602), .Q(
        \gbuff[30][0] ) );
  DFFRX1 \gbuff_reg[26][31]  ( .D(n1955), .CK(clk), .RN(n1593), .Q(
        \gbuff[26][31] ) );
  DFFRX1 \gbuff_reg[26][30]  ( .D(n1956), .CK(clk), .RN(n1593), .Q(
        \gbuff[26][30] ) );
  DFFRX1 \gbuff_reg[26][29]  ( .D(n1957), .CK(clk), .RN(n1593), .Q(
        \gbuff[26][29] ) );
  DFFRX1 \gbuff_reg[26][28]  ( .D(n1958), .CK(clk), .RN(n1593), .Q(
        \gbuff[26][28] ) );
  DFFRX1 \gbuff_reg[26][27]  ( .D(n1959), .CK(clk), .RN(n1593), .Q(
        \gbuff[26][27] ) );
  DFFRX1 \gbuff_reg[26][26]  ( .D(n1960), .CK(clk), .RN(n1593), .Q(
        \gbuff[26][26] ) );
  DFFRX1 \gbuff_reg[26][25]  ( .D(n1961), .CK(clk), .RN(n1593), .Q(
        \gbuff[26][25] ) );
  DFFRX1 \gbuff_reg[26][24]  ( .D(n1962), .CK(clk), .RN(n1593), .Q(
        \gbuff[26][24] ) );
  DFFRX1 \gbuff_reg[26][23]  ( .D(n1963), .CK(clk), .RN(n1593), .Q(
        \gbuff[26][23] ) );
  DFFRX1 \gbuff_reg[26][22]  ( .D(n1964), .CK(clk), .RN(n1593), .Q(
        \gbuff[26][22] ) );
  DFFRX1 \gbuff_reg[26][21]  ( .D(n1965), .CK(clk), .RN(n1593), .Q(
        \gbuff[26][21] ) );
  DFFRX1 \gbuff_reg[26][20]  ( .D(n1966), .CK(clk), .RN(n1593), .Q(
        \gbuff[26][20] ) );
  DFFRX1 \gbuff_reg[26][19]  ( .D(n1967), .CK(clk), .RN(n1592), .Q(
        \gbuff[26][19] ) );
  DFFRX1 \gbuff_reg[26][18]  ( .D(n1968), .CK(clk), .RN(n1592), .Q(
        \gbuff[26][18] ) );
  DFFRX1 \gbuff_reg[26][17]  ( .D(n1969), .CK(clk), .RN(n1592), .Q(
        \gbuff[26][17] ) );
  DFFRX1 \gbuff_reg[26][16]  ( .D(n1970), .CK(clk), .RN(n1592), .Q(
        \gbuff[26][16] ) );
  DFFRX1 \gbuff_reg[26][15]  ( .D(n1971), .CK(clk), .RN(n1592), .Q(
        \gbuff[26][15] ) );
  DFFRX1 \gbuff_reg[26][14]  ( .D(n1972), .CK(clk), .RN(n1592), .Q(
        \gbuff[26][14] ) );
  DFFRX1 \gbuff_reg[26][13]  ( .D(n1973), .CK(clk), .RN(n1592), .Q(
        \gbuff[26][13] ) );
  DFFRX1 \gbuff_reg[26][12]  ( .D(n1974), .CK(clk), .RN(n1592), .Q(
        \gbuff[26][12] ) );
  DFFRX1 \gbuff_reg[26][11]  ( .D(n1975), .CK(clk), .RN(n1592), .Q(
        \gbuff[26][11] ) );
  DFFRX1 \gbuff_reg[26][10]  ( .D(n1976), .CK(clk), .RN(n1592), .Q(
        \gbuff[26][10] ) );
  DFFRX1 \gbuff_reg[26][9]  ( .D(n1977), .CK(clk), .RN(n1592), .Q(
        \gbuff[26][9] ) );
  DFFRX1 \gbuff_reg[26][8]  ( .D(n1978), .CK(clk), .RN(n1592), .Q(
        \gbuff[26][8] ) );
  DFFRX1 \gbuff_reg[26][7]  ( .D(n1979), .CK(clk), .RN(n1591), .Q(
        \gbuff[26][7] ) );
  DFFRX1 \gbuff_reg[26][6]  ( .D(n1980), .CK(clk), .RN(n1591), .Q(
        \gbuff[26][6] ) );
  DFFRX1 \gbuff_reg[26][5]  ( .D(n1981), .CK(clk), .RN(n1591), .Q(
        \gbuff[26][5] ) );
  DFFRX1 \gbuff_reg[26][4]  ( .D(n1982), .CK(clk), .RN(n1591), .Q(
        \gbuff[26][4] ) );
  DFFRX1 \gbuff_reg[26][3]  ( .D(n1983), .CK(clk), .RN(n1591), .Q(
        \gbuff[26][3] ) );
  DFFRX1 \gbuff_reg[26][2]  ( .D(n1984), .CK(clk), .RN(n1591), .Q(
        \gbuff[26][2] ) );
  DFFRX1 \gbuff_reg[26][1]  ( .D(n1985), .CK(clk), .RN(n1591), .Q(
        \gbuff[26][1] ) );
  DFFRX1 \gbuff_reg[26][0]  ( .D(n1986), .CK(clk), .RN(n1591), .Q(
        \gbuff[26][0] ) );
  DFFRX1 \gbuff_reg[22][31]  ( .D(n2083), .CK(clk), .RN(n1583), .Q(
        \gbuff[22][31] ) );
  DFFRX1 \gbuff_reg[22][30]  ( .D(n2084), .CK(clk), .RN(n1583), .Q(
        \gbuff[22][30] ) );
  DFFRX1 \gbuff_reg[22][29]  ( .D(n2085), .CK(clk), .RN(n1583), .Q(
        \gbuff[22][29] ) );
  DFFRX1 \gbuff_reg[22][28]  ( .D(n2086), .CK(clk), .RN(n1583), .Q(
        \gbuff[22][28] ) );
  DFFRX1 \gbuff_reg[22][27]  ( .D(n2087), .CK(clk), .RN(n1582), .Q(
        \gbuff[22][27] ) );
  DFFRX1 \gbuff_reg[22][26]  ( .D(n2088), .CK(clk), .RN(n1582), .Q(
        \gbuff[22][26] ) );
  DFFRX1 \gbuff_reg[22][25]  ( .D(n2089), .CK(clk), .RN(n1582), .Q(
        \gbuff[22][25] ) );
  DFFRX1 \gbuff_reg[22][24]  ( .D(n2090), .CK(clk), .RN(n1582), .Q(
        \gbuff[22][24] ) );
  DFFRX1 \gbuff_reg[22][23]  ( .D(n2091), .CK(clk), .RN(n1582), .Q(
        \gbuff[22][23] ) );
  DFFRX1 \gbuff_reg[22][22]  ( .D(n2092), .CK(clk), .RN(n1582), .Q(
        \gbuff[22][22] ) );
  DFFRX1 \gbuff_reg[22][21]  ( .D(n2093), .CK(clk), .RN(n1582), .Q(
        \gbuff[22][21] ) );
  DFFRX1 \gbuff_reg[22][20]  ( .D(n2094), .CK(clk), .RN(n1582), .Q(
        \gbuff[22][20] ) );
  DFFRX1 \gbuff_reg[22][19]  ( .D(n2095), .CK(clk), .RN(n1582), .Q(
        \gbuff[22][19] ) );
  DFFRX1 \gbuff_reg[22][18]  ( .D(n2096), .CK(clk), .RN(n1582), .Q(
        \gbuff[22][18] ) );
  DFFRX1 \gbuff_reg[22][17]  ( .D(n2097), .CK(clk), .RN(n1582), .Q(
        \gbuff[22][17] ) );
  DFFRX1 \gbuff_reg[22][16]  ( .D(n2098), .CK(clk), .RN(n1582), .Q(
        \gbuff[22][16] ) );
  DFFRX1 \gbuff_reg[22][15]  ( .D(n2099), .CK(clk), .RN(n1581), .Q(
        \gbuff[22][15] ) );
  DFFRX1 \gbuff_reg[22][14]  ( .D(n2100), .CK(clk), .RN(n1581), .Q(
        \gbuff[22][14] ) );
  DFFRX1 \gbuff_reg[22][13]  ( .D(n2101), .CK(clk), .RN(n1581), .Q(
        \gbuff[22][13] ) );
  DFFRX1 \gbuff_reg[22][12]  ( .D(n2102), .CK(clk), .RN(n1581), .Q(
        \gbuff[22][12] ) );
  DFFRX1 \gbuff_reg[22][11]  ( .D(n2103), .CK(clk), .RN(n1581), .Q(
        \gbuff[22][11] ) );
  DFFRX1 \gbuff_reg[22][10]  ( .D(n2104), .CK(clk), .RN(n1581), .Q(
        \gbuff[22][10] ) );
  DFFRX1 \gbuff_reg[22][9]  ( .D(n2105), .CK(clk), .RN(n1581), .Q(
        \gbuff[22][9] ) );
  DFFRX1 \gbuff_reg[22][8]  ( .D(n2106), .CK(clk), .RN(n1581), .Q(
        \gbuff[22][8] ) );
  DFFRX1 \gbuff_reg[22][7]  ( .D(n2107), .CK(clk), .RN(n1581), .Q(
        \gbuff[22][7] ) );
  DFFRX1 \gbuff_reg[22][6]  ( .D(n2108), .CK(clk), .RN(n1581), .Q(
        \gbuff[22][6] ) );
  DFFRX1 \gbuff_reg[22][5]  ( .D(n2109), .CK(clk), .RN(n1581), .Q(
        \gbuff[22][5] ) );
  DFFRX1 \gbuff_reg[22][4]  ( .D(n2110), .CK(clk), .RN(n1581), .Q(
        \gbuff[22][4] ) );
  DFFRX1 \gbuff_reg[22][3]  ( .D(n2111), .CK(clk), .RN(n1580), .Q(
        \gbuff[22][3] ) );
  DFFRX1 \gbuff_reg[22][2]  ( .D(n2112), .CK(clk), .RN(n1580), .Q(
        \gbuff[22][2] ) );
  DFFRX1 \gbuff_reg[22][1]  ( .D(n2113), .CK(clk), .RN(n1580), .Q(
        \gbuff[22][1] ) );
  DFFRX1 \gbuff_reg[22][0]  ( .D(n2114), .CK(clk), .RN(n1580), .Q(
        \gbuff[22][0] ) );
  DFFRX1 \gbuff_reg[18][31]  ( .D(n2211), .CK(clk), .RN(n1572), .Q(
        \gbuff[18][31] ) );
  DFFRX1 \gbuff_reg[18][30]  ( .D(n2212), .CK(clk), .RN(n1572), .Q(
        \gbuff[18][30] ) );
  DFFRX1 \gbuff_reg[18][29]  ( .D(n2213), .CK(clk), .RN(n1572), .Q(
        \gbuff[18][29] ) );
  DFFRX1 \gbuff_reg[18][28]  ( .D(n2214), .CK(clk), .RN(n1572), .Q(
        \gbuff[18][28] ) );
  DFFRX1 \gbuff_reg[18][27]  ( .D(n2215), .CK(clk), .RN(n1572), .Q(
        \gbuff[18][27] ) );
  DFFRX1 \gbuff_reg[18][26]  ( .D(n2216), .CK(clk), .RN(n1572), .Q(
        \gbuff[18][26] ) );
  DFFRX1 \gbuff_reg[18][25]  ( .D(n2217), .CK(clk), .RN(n1572), .Q(
        \gbuff[18][25] ) );
  DFFRX1 \gbuff_reg[18][24]  ( .D(n2218), .CK(clk), .RN(n1572), .Q(
        \gbuff[18][24] ) );
  DFFRX1 \gbuff_reg[18][23]  ( .D(n2219), .CK(clk), .RN(n1571), .Q(
        \gbuff[18][23] ) );
  DFFRX1 \gbuff_reg[18][22]  ( .D(n2220), .CK(clk), .RN(n1571), .Q(
        \gbuff[18][22] ) );
  DFFRX1 \gbuff_reg[18][21]  ( .D(n2221), .CK(clk), .RN(n1571), .Q(
        \gbuff[18][21] ) );
  DFFRX1 \gbuff_reg[18][20]  ( .D(n2222), .CK(clk), .RN(n1571), .Q(
        \gbuff[18][20] ) );
  DFFRX1 \gbuff_reg[18][19]  ( .D(n2223), .CK(clk), .RN(n1571), .Q(
        \gbuff[18][19] ) );
  DFFRX1 \gbuff_reg[18][18]  ( .D(n2224), .CK(clk), .RN(n1571), .Q(
        \gbuff[18][18] ) );
  DFFRX1 \gbuff_reg[18][17]  ( .D(n2225), .CK(clk), .RN(n1571), .Q(
        \gbuff[18][17] ) );
  DFFRX1 \gbuff_reg[18][16]  ( .D(n2226), .CK(clk), .RN(n1571), .Q(
        \gbuff[18][16] ) );
  DFFRX1 \gbuff_reg[18][15]  ( .D(n2227), .CK(clk), .RN(n1571), .Q(
        \gbuff[18][15] ) );
  DFFRX1 \gbuff_reg[18][14]  ( .D(n2228), .CK(clk), .RN(n1571), .Q(
        \gbuff[18][14] ) );
  DFFRX1 \gbuff_reg[18][13]  ( .D(n2229), .CK(clk), .RN(n1571), .Q(
        \gbuff[18][13] ) );
  DFFRX1 \gbuff_reg[18][12]  ( .D(n2230), .CK(clk), .RN(n1571), .Q(
        \gbuff[18][12] ) );
  DFFRX1 \gbuff_reg[18][11]  ( .D(n2231), .CK(clk), .RN(n1570), .Q(
        \gbuff[18][11] ) );
  DFFRX1 \gbuff_reg[18][10]  ( .D(n2232), .CK(clk), .RN(n1570), .Q(
        \gbuff[18][10] ) );
  DFFRX1 \gbuff_reg[18][9]  ( .D(n2233), .CK(clk), .RN(n1570), .Q(
        \gbuff[18][9] ) );
  DFFRX1 \gbuff_reg[18][8]  ( .D(n2234), .CK(clk), .RN(n1570), .Q(
        \gbuff[18][8] ) );
  DFFRX1 \gbuff_reg[18][7]  ( .D(n2235), .CK(clk), .RN(n1570), .Q(
        \gbuff[18][7] ) );
  DFFRX1 \gbuff_reg[18][6]  ( .D(n2236), .CK(clk), .RN(n1570), .Q(
        \gbuff[18][6] ) );
  DFFRX1 \gbuff_reg[18][5]  ( .D(n2237), .CK(clk), .RN(n1570), .Q(
        \gbuff[18][5] ) );
  DFFRX1 \gbuff_reg[18][4]  ( .D(n2238), .CK(clk), .RN(n1570), .Q(
        \gbuff[18][4] ) );
  DFFRX1 \gbuff_reg[18][3]  ( .D(n2239), .CK(clk), .RN(n1570), .Q(
        \gbuff[18][3] ) );
  DFFRX1 \gbuff_reg[18][2]  ( .D(n2240), .CK(clk), .RN(n1570), .Q(
        \gbuff[18][2] ) );
  DFFRX1 \gbuff_reg[18][1]  ( .D(n2241), .CK(clk), .RN(n1570), .Q(
        \gbuff[18][1] ) );
  DFFRX1 \gbuff_reg[18][0]  ( .D(n2242), .CK(clk), .RN(n1570), .Q(
        \gbuff[18][0] ) );
  DFFRX1 \gbuff_reg[14][31]  ( .D(n2339), .CK(clk), .RN(n1561), .Q(
        \gbuff[14][31] ) );
  DFFRX1 \gbuff_reg[14][30]  ( .D(n2340), .CK(clk), .RN(n1561), .Q(
        \gbuff[14][30] ) );
  DFFRX1 \gbuff_reg[14][29]  ( .D(n2341), .CK(clk), .RN(n1561), .Q(
        \gbuff[14][29] ) );
  DFFRX1 \gbuff_reg[14][28]  ( .D(n2342), .CK(clk), .RN(n1561), .Q(
        \gbuff[14][28] ) );
  DFFRX1 \gbuff_reg[14][27]  ( .D(n2343), .CK(clk), .RN(n1561), .Q(
        \gbuff[14][27] ) );
  DFFRX1 \gbuff_reg[14][26]  ( .D(n2344), .CK(clk), .RN(n1561), .Q(
        \gbuff[14][26] ) );
  DFFRX1 \gbuff_reg[14][25]  ( .D(n2345), .CK(clk), .RN(n1561), .Q(
        \gbuff[14][25] ) );
  DFFRX1 \gbuff_reg[14][24]  ( .D(n2346), .CK(clk), .RN(n1561), .Q(
        \gbuff[14][24] ) );
  DFFRX1 \gbuff_reg[14][23]  ( .D(n2347), .CK(clk), .RN(n1561), .Q(
        \gbuff[14][23] ) );
  DFFRX1 \gbuff_reg[14][22]  ( .D(n2348), .CK(clk), .RN(n1561), .Q(
        \gbuff[14][22] ) );
  DFFRX1 \gbuff_reg[14][21]  ( .D(n2349), .CK(clk), .RN(n1561), .Q(
        \gbuff[14][21] ) );
  DFFRX1 \gbuff_reg[14][20]  ( .D(n2350), .CK(clk), .RN(n1561), .Q(
        \gbuff[14][20] ) );
  DFFRX1 \gbuff_reg[14][19]  ( .D(n2351), .CK(clk), .RN(n1560), .Q(
        \gbuff[14][19] ) );
  DFFRX1 \gbuff_reg[14][18]  ( .D(n2352), .CK(clk), .RN(n1560), .Q(
        \gbuff[14][18] ) );
  DFFRX1 \gbuff_reg[14][17]  ( .D(n2353), .CK(clk), .RN(n1560), .Q(
        \gbuff[14][17] ) );
  DFFRX1 \gbuff_reg[14][16]  ( .D(n2354), .CK(clk), .RN(n1560), .Q(
        \gbuff[14][16] ) );
  DFFRX1 \gbuff_reg[14][15]  ( .D(n2355), .CK(clk), .RN(n1560), .Q(
        \gbuff[14][15] ) );
  DFFRX1 \gbuff_reg[14][14]  ( .D(n2356), .CK(clk), .RN(n1560), .Q(
        \gbuff[14][14] ) );
  DFFRX1 \gbuff_reg[14][13]  ( .D(n2357), .CK(clk), .RN(n1560), .Q(
        \gbuff[14][13] ) );
  DFFRX1 \gbuff_reg[14][12]  ( .D(n2358), .CK(clk), .RN(n1560), .Q(
        \gbuff[14][12] ) );
  DFFRX1 \gbuff_reg[14][11]  ( .D(n2359), .CK(clk), .RN(n1560), .Q(
        \gbuff[14][11] ) );
  DFFRX1 \gbuff_reg[14][10]  ( .D(n2360), .CK(clk), .RN(n1560), .Q(
        \gbuff[14][10] ) );
  DFFRX1 \gbuff_reg[14][9]  ( .D(n2361), .CK(clk), .RN(n1560), .Q(
        \gbuff[14][9] ) );
  DFFRX1 \gbuff_reg[14][8]  ( .D(n2362), .CK(clk), .RN(n1560), .Q(
        \gbuff[14][8] ) );
  DFFRX1 \gbuff_reg[14][7]  ( .D(n2363), .CK(clk), .RN(n1559), .Q(
        \gbuff[14][7] ) );
  DFFRX1 \gbuff_reg[14][6]  ( .D(n2364), .CK(clk), .RN(n1559), .Q(
        \gbuff[14][6] ) );
  DFFRX1 \gbuff_reg[14][5]  ( .D(n2365), .CK(clk), .RN(n1559), .Q(
        \gbuff[14][5] ) );
  DFFRX1 \gbuff_reg[14][4]  ( .D(n2366), .CK(clk), .RN(n1559), .Q(
        \gbuff[14][4] ) );
  DFFRX1 \gbuff_reg[14][3]  ( .D(n2367), .CK(clk), .RN(n1559), .Q(
        \gbuff[14][3] ) );
  DFFRX1 \gbuff_reg[14][2]  ( .D(n2368), .CK(clk), .RN(n1559), .Q(
        \gbuff[14][2] ) );
  DFFRX1 \gbuff_reg[14][1]  ( .D(n2369), .CK(clk), .RN(n1559), .Q(
        \gbuff[14][1] ) );
  DFFRX1 \gbuff_reg[14][0]  ( .D(n2370), .CK(clk), .RN(n1559), .Q(
        \gbuff[14][0] ) );
  DFFRX1 \gbuff_reg[10][31]  ( .D(n2467), .CK(clk), .RN(n1551), .Q(
        \gbuff[10][31] ) );
  DFFRX1 \gbuff_reg[10][30]  ( .D(n2468), .CK(clk), .RN(n1551), .Q(
        \gbuff[10][30] ) );
  DFFRX1 \gbuff_reg[10][29]  ( .D(n2469), .CK(clk), .RN(n1551), .Q(
        \gbuff[10][29] ) );
  DFFRX1 \gbuff_reg[10][28]  ( .D(n2470), .CK(clk), .RN(n1551), .Q(
        \gbuff[10][28] ) );
  DFFRX1 \gbuff_reg[10][27]  ( .D(n2471), .CK(clk), .RN(n1550), .Q(
        \gbuff[10][27] ) );
  DFFRX1 \gbuff_reg[10][26]  ( .D(n2472), .CK(clk), .RN(n1550), .Q(
        \gbuff[10][26] ) );
  DFFRX1 \gbuff_reg[10][25]  ( .D(n2473), .CK(clk), .RN(n1550), .Q(
        \gbuff[10][25] ) );
  DFFRX1 \gbuff_reg[10][24]  ( .D(n2474), .CK(clk), .RN(n1550), .Q(
        \gbuff[10][24] ) );
  DFFRX1 \gbuff_reg[10][23]  ( .D(n2475), .CK(clk), .RN(n1550), .Q(
        \gbuff[10][23] ) );
  DFFRX1 \gbuff_reg[10][22]  ( .D(n2476), .CK(clk), .RN(n1550), .Q(
        \gbuff[10][22] ) );
  DFFRX1 \gbuff_reg[10][21]  ( .D(n2477), .CK(clk), .RN(n1550), .Q(
        \gbuff[10][21] ) );
  DFFRX1 \gbuff_reg[10][20]  ( .D(n2478), .CK(clk), .RN(n1550), .Q(
        \gbuff[10][20] ) );
  DFFRX1 \gbuff_reg[10][19]  ( .D(n2479), .CK(clk), .RN(n1550), .Q(
        \gbuff[10][19] ) );
  DFFRX1 \gbuff_reg[10][18]  ( .D(n2480), .CK(clk), .RN(n1550), .Q(
        \gbuff[10][18] ) );
  DFFRX1 \gbuff_reg[10][17]  ( .D(n2481), .CK(clk), .RN(n1550), .Q(
        \gbuff[10][17] ) );
  DFFRX1 \gbuff_reg[10][16]  ( .D(n2482), .CK(clk), .RN(n1550), .Q(
        \gbuff[10][16] ) );
  DFFRX1 \gbuff_reg[10][15]  ( .D(n2483), .CK(clk), .RN(n1549), .Q(
        \gbuff[10][15] ) );
  DFFRX1 \gbuff_reg[10][14]  ( .D(n2484), .CK(clk), .RN(n1549), .Q(
        \gbuff[10][14] ) );
  DFFRX1 \gbuff_reg[10][13]  ( .D(n2485), .CK(clk), .RN(n1549), .Q(
        \gbuff[10][13] ) );
  DFFRX1 \gbuff_reg[10][12]  ( .D(n2486), .CK(clk), .RN(n1549), .Q(
        \gbuff[10][12] ) );
  DFFRX1 \gbuff_reg[10][11]  ( .D(n2487), .CK(clk), .RN(n1549), .Q(
        \gbuff[10][11] ) );
  DFFRX1 \gbuff_reg[10][10]  ( .D(n2488), .CK(clk), .RN(n1549), .Q(
        \gbuff[10][10] ) );
  DFFRX1 \gbuff_reg[10][9]  ( .D(n2489), .CK(clk), .RN(n1549), .Q(
        \gbuff[10][9] ) );
  DFFRX1 \gbuff_reg[10][8]  ( .D(n2490), .CK(clk), .RN(n1549), .Q(
        \gbuff[10][8] ) );
  DFFRX1 \gbuff_reg[10][7]  ( .D(n2491), .CK(clk), .RN(n1549), .Q(
        \gbuff[10][7] ) );
  DFFRX1 \gbuff_reg[10][6]  ( .D(n2492), .CK(clk), .RN(n1549), .Q(
        \gbuff[10][6] ) );
  DFFRX1 \gbuff_reg[10][5]  ( .D(n2493), .CK(clk), .RN(n1549), .Q(
        \gbuff[10][5] ) );
  DFFRX1 \gbuff_reg[10][4]  ( .D(n2494), .CK(clk), .RN(n1549), .Q(
        \gbuff[10][4] ) );
  DFFRX1 \gbuff_reg[10][3]  ( .D(n2495), .CK(clk), .RN(n1548), .Q(
        \gbuff[10][3] ) );
  DFFRX1 \gbuff_reg[10][2]  ( .D(n2496), .CK(clk), .RN(n1548), .Q(
        \gbuff[10][2] ) );
  DFFRX1 \gbuff_reg[10][1]  ( .D(n2497), .CK(clk), .RN(n1548), .Q(
        \gbuff[10][1] ) );
  DFFRX1 \gbuff_reg[10][0]  ( .D(n2498), .CK(clk), .RN(n1548), .Q(
        \gbuff[10][0] ) );
  DFFRX1 \gbuff_reg[6][31]  ( .D(n2595), .CK(clk), .RN(n1540), .Q(
        \gbuff[6][31] ) );
  DFFRX1 \gbuff_reg[6][30]  ( .D(n2596), .CK(clk), .RN(n1540), .Q(
        \gbuff[6][30] ) );
  DFFRX1 \gbuff_reg[6][29]  ( .D(n2597), .CK(clk), .RN(n1540), .Q(
        \gbuff[6][29] ) );
  DFFRX1 \gbuff_reg[6][28]  ( .D(n2598), .CK(clk), .RN(n1540), .Q(
        \gbuff[6][28] ) );
  DFFRX1 \gbuff_reg[6][27]  ( .D(n2599), .CK(clk), .RN(n1540), .Q(
        \gbuff[6][27] ) );
  DFFRX1 \gbuff_reg[6][26]  ( .D(n2600), .CK(clk), .RN(n1540), .Q(
        \gbuff[6][26] ) );
  DFFRX1 \gbuff_reg[6][25]  ( .D(n2601), .CK(clk), .RN(n1540), .Q(
        \gbuff[6][25] ) );
  DFFRX1 \gbuff_reg[6][24]  ( .D(n2602), .CK(clk), .RN(n1540), .Q(
        \gbuff[6][24] ) );
  DFFRX1 \gbuff_reg[6][23]  ( .D(n2603), .CK(clk), .RN(n1539), .Q(
        \gbuff[6][23] ) );
  DFFRX1 \gbuff_reg[6][22]  ( .D(n2604), .CK(clk), .RN(n1539), .Q(
        \gbuff[6][22] ) );
  DFFRX1 \gbuff_reg[6][21]  ( .D(n2605), .CK(clk), .RN(n1539), .Q(
        \gbuff[6][21] ) );
  DFFRX1 \gbuff_reg[6][20]  ( .D(n2606), .CK(clk), .RN(n1539), .Q(
        \gbuff[6][20] ) );
  DFFRX1 \gbuff_reg[6][19]  ( .D(n2607), .CK(clk), .RN(n1539), .Q(
        \gbuff[6][19] ) );
  DFFRX1 \gbuff_reg[6][18]  ( .D(n2608), .CK(clk), .RN(n1539), .Q(
        \gbuff[6][18] ) );
  DFFRX1 \gbuff_reg[6][17]  ( .D(n2609), .CK(clk), .RN(n1539), .Q(
        \gbuff[6][17] ) );
  DFFRX1 \gbuff_reg[6][16]  ( .D(n2610), .CK(clk), .RN(n1539), .Q(
        \gbuff[6][16] ) );
  DFFRX1 \gbuff_reg[6][15]  ( .D(n2611), .CK(clk), .RN(n1539), .Q(
        \gbuff[6][15] ) );
  DFFRX1 \gbuff_reg[6][14]  ( .D(n2612), .CK(clk), .RN(n1539), .Q(
        \gbuff[6][14] ) );
  DFFRX1 \gbuff_reg[6][13]  ( .D(n2613), .CK(clk), .RN(n1539), .Q(
        \gbuff[6][13] ) );
  DFFRX1 \gbuff_reg[6][12]  ( .D(n2614), .CK(clk), .RN(n1539), .Q(
        \gbuff[6][12] ) );
  DFFRX1 \gbuff_reg[6][11]  ( .D(n2615), .CK(clk), .RN(n1538), .Q(
        \gbuff[6][11] ) );
  DFFRX1 \gbuff_reg[6][10]  ( .D(n2616), .CK(clk), .RN(n1538), .Q(
        \gbuff[6][10] ) );
  DFFRX1 \gbuff_reg[6][9]  ( .D(n2617), .CK(clk), .RN(n1538), .Q(\gbuff[6][9] ) );
  DFFRX1 \gbuff_reg[6][8]  ( .D(n2618), .CK(clk), .RN(n1538), .Q(\gbuff[6][8] ) );
  DFFRX1 \gbuff_reg[6][7]  ( .D(n2619), .CK(clk), .RN(n1538), .Q(\gbuff[6][7] ) );
  DFFRX1 \gbuff_reg[6][6]  ( .D(n2620), .CK(clk), .RN(n1538), .Q(\gbuff[6][6] ) );
  DFFRX1 \gbuff_reg[6][5]  ( .D(n2621), .CK(clk), .RN(n1538), .Q(\gbuff[6][5] ) );
  DFFRX1 \gbuff_reg[6][4]  ( .D(n2622), .CK(clk), .RN(n1538), .Q(\gbuff[6][4] ) );
  DFFRX1 \gbuff_reg[6][3]  ( .D(n2623), .CK(clk), .RN(n1538), .Q(\gbuff[6][3] ) );
  DFFRX1 \gbuff_reg[6][2]  ( .D(n2624), .CK(clk), .RN(n1538), .Q(\gbuff[6][2] ) );
  DFFRX1 \gbuff_reg[6][1]  ( .D(n2625), .CK(clk), .RN(n1538), .Q(\gbuff[6][1] ) );
  DFFRX1 \gbuff_reg[6][0]  ( .D(n2626), .CK(clk), .RN(n1538), .Q(\gbuff[6][0] ) );
  DFFRX1 \gbuff_reg[2][31]  ( .D(n2723), .CK(clk), .RN(n1529), .Q(
        \gbuff[2][31] ) );
  DFFRX1 \gbuff_reg[2][30]  ( .D(n2724), .CK(clk), .RN(n1529), .Q(
        \gbuff[2][30] ) );
  DFFRX1 \gbuff_reg[2][29]  ( .D(n2725), .CK(clk), .RN(n1529), .Q(
        \gbuff[2][29] ) );
  DFFRX1 \gbuff_reg[2][28]  ( .D(n2726), .CK(clk), .RN(n1529), .Q(
        \gbuff[2][28] ) );
  DFFRX1 \gbuff_reg[2][27]  ( .D(n2727), .CK(clk), .RN(n1529), .Q(
        \gbuff[2][27] ) );
  DFFRX1 \gbuff_reg[2][26]  ( .D(n2728), .CK(clk), .RN(n1529), .Q(
        \gbuff[2][26] ) );
  DFFRX1 \gbuff_reg[2][25]  ( .D(n2729), .CK(clk), .RN(n1529), .Q(
        \gbuff[2][25] ) );
  DFFRX1 \gbuff_reg[2][24]  ( .D(n2730), .CK(clk), .RN(n1529), .Q(
        \gbuff[2][24] ) );
  DFFRX1 \gbuff_reg[2][23]  ( .D(n2731), .CK(clk), .RN(n1529), .Q(
        \gbuff[2][23] ) );
  DFFRX1 \gbuff_reg[2][22]  ( .D(n2732), .CK(clk), .RN(n1529), .Q(
        \gbuff[2][22] ) );
  DFFRX1 \gbuff_reg[2][21]  ( .D(n2733), .CK(clk), .RN(n1529), .Q(
        \gbuff[2][21] ) );
  DFFRX1 \gbuff_reg[2][20]  ( .D(n2734), .CK(clk), .RN(n1529), .Q(
        \gbuff[2][20] ) );
  DFFRX1 \gbuff_reg[2][19]  ( .D(n2735), .CK(clk), .RN(n1528), .Q(
        \gbuff[2][19] ) );
  DFFRX1 \gbuff_reg[2][18]  ( .D(n2736), .CK(clk), .RN(n1528), .Q(
        \gbuff[2][18] ) );
  DFFRX1 \gbuff_reg[2][17]  ( .D(n2737), .CK(clk), .RN(n1528), .Q(
        \gbuff[2][17] ) );
  DFFRX1 \gbuff_reg[2][16]  ( .D(n2738), .CK(clk), .RN(n1528), .Q(
        \gbuff[2][16] ) );
  DFFRX1 \gbuff_reg[2][15]  ( .D(n2739), .CK(clk), .RN(n1528), .Q(
        \gbuff[2][15] ) );
  DFFRX1 \gbuff_reg[2][14]  ( .D(n2740), .CK(clk), .RN(n1528), .Q(
        \gbuff[2][14] ) );
  DFFRX1 \gbuff_reg[2][13]  ( .D(n2741), .CK(clk), .RN(n1528), .Q(
        \gbuff[2][13] ) );
  DFFRX1 \gbuff_reg[2][12]  ( .D(n2742), .CK(clk), .RN(n1528), .Q(
        \gbuff[2][12] ) );
  DFFRX1 \gbuff_reg[2][11]  ( .D(n2743), .CK(clk), .RN(n1528), .Q(
        \gbuff[2][11] ) );
  DFFRX1 \gbuff_reg[2][10]  ( .D(n2744), .CK(clk), .RN(n1528), .Q(
        \gbuff[2][10] ) );
  DFFRX1 \gbuff_reg[2][9]  ( .D(n2745), .CK(clk), .RN(n1528), .Q(\gbuff[2][9] ) );
  DFFRX1 \gbuff_reg[2][8]  ( .D(n2746), .CK(clk), .RN(n1528), .Q(\gbuff[2][8] ) );
  DFFRX1 \gbuff_reg[2][7]  ( .D(n2747), .CK(clk), .RN(n1527), .Q(\gbuff[2][7] ) );
  DFFRX1 \gbuff_reg[2][6]  ( .D(n2748), .CK(clk), .RN(n1527), .Q(\gbuff[2][6] ) );
  DFFRX1 \gbuff_reg[2][5]  ( .D(n2749), .CK(clk), .RN(n1527), .Q(\gbuff[2][5] ) );
  DFFRX1 \gbuff_reg[2][4]  ( .D(n2750), .CK(clk), .RN(n1527), .Q(\gbuff[2][4] ) );
  DFFRX1 \gbuff_reg[2][3]  ( .D(n2751), .CK(clk), .RN(n1527), .Q(\gbuff[2][3] ) );
  DFFRX1 \gbuff_reg[2][2]  ( .D(n2752), .CK(clk), .RN(n1527), .Q(\gbuff[2][2] ) );
  DFFRX1 \gbuff_reg[2][1]  ( .D(n2753), .CK(clk), .RN(n1527), .Q(\gbuff[2][1] ) );
  DFFRX1 \gbuff_reg[2][0]  ( .D(n2754), .CK(clk), .RN(n1527), .Q(\gbuff[2][0] ) );
  EDFFTRX2 \data_out_reg[19]  ( .RN(1'b1), .D(N28), .E(N81), .CK(clk), .Q(
        data_out[19]) );
  EDFFTRX2 \data_out_reg[18]  ( .RN(1'b1), .D(N29), .E(N81), .CK(clk), .Q(
        data_out[18]) );
  EDFFTRX2 \data_out_reg[17]  ( .RN(1'b1), .D(N30), .E(N81), .CK(clk), .Q(
        data_out[17]) );
  EDFFTRX2 \data_out_reg[16]  ( .RN(1'b1), .D(N31), .E(N81), .CK(clk), .Q(
        data_out[16]) );
  EDFFTRX2 \data_out_reg[31]  ( .RN(1'b1), .D(N16), .E(N81), .CK(clk), .Q(
        data_out[31]) );
  EDFFTRX2 \data_out_reg[30]  ( .RN(1'b1), .D(N17), .E(N81), .CK(clk), .Q(
        data_out[30]) );
  EDFFTRX2 \data_out_reg[29]  ( .RN(1'b1), .D(N18), .E(N81), .CK(clk), .Q(
        data_out[29]) );
  EDFFTRX2 \data_out_reg[28]  ( .RN(1'b1), .D(N19), .E(N81), .CK(clk), .Q(
        data_out[28]) );
  EDFFTRX2 \data_out_reg[27]  ( .RN(1'b1), .D(N20), .E(N81), .CK(clk), .Q(
        data_out[27]) );
  EDFFTRX2 \data_out_reg[26]  ( .RN(1'b1), .D(N21), .E(N81), .CK(clk), .Q(
        data_out[26]) );
  EDFFTRX2 \data_out_reg[25]  ( .RN(1'b1), .D(N22), .E(N81), .CK(clk), .Q(
        data_out[25]) );
  EDFFTRX2 \data_out_reg[24]  ( .RN(1'b1), .D(N23), .E(N81), .CK(clk), .Q(
        data_out[24]) );
  EDFFTRX2 \data_out_reg[23]  ( .RN(1'b1), .D(N24), .E(N81), .CK(clk), .Q(
        data_out[23]) );
  EDFFTRX2 \data_out_reg[22]  ( .RN(1'b1), .D(N25), .E(N81), .CK(clk), .Q(
        data_out[22]) );
  EDFFTRX2 \data_out_reg[21]  ( .RN(1'b1), .D(N26), .E(N81), .CK(clk), .Q(
        data_out[21]) );
  EDFFTRX2 \data_out_reg[20]  ( .RN(1'b1), .D(N27), .E(N81), .CK(clk), .Q(
        data_out[20]) );
  EDFFX2 \data_out_reg[15]  ( .D(N32), .E(N81), .CK(clk), .Q(data_out[15]) );
  EDFFX2 \data_out_reg[14]  ( .D(N33), .E(N81), .CK(clk), .Q(data_out[14]) );
  EDFFX2 \data_out_reg[13]  ( .D(N34), .E(N81), .CK(clk), .Q(data_out[13]) );
  EDFFX2 \data_out_reg[12]  ( .D(N35), .E(n1755), .CK(clk), .Q(data_out[12])
         );
  EDFFX2 \data_out_reg[11]  ( .D(N36), .E(n1755), .CK(clk), .Q(data_out[11])
         );
  EDFFX2 \data_out_reg[10]  ( .D(N37), .E(n1755), .CK(clk), .Q(data_out[10])
         );
  EDFFX2 \data_out_reg[9]  ( .D(N38), .E(n1755), .CK(clk), .Q(data_out[9]) );
  EDFFX2 \data_out_reg[8]  ( .D(N39), .E(n1755), .CK(clk), .Q(data_out[8]) );
  EDFFX2 \data_out_reg[7]  ( .D(N40), .E(n1755), .CK(clk), .Q(data_out[7]) );
  EDFFX2 \data_out_reg[6]  ( .D(N41), .E(n1755), .CK(clk), .Q(data_out[6]) );
  EDFFX2 \data_out_reg[5]  ( .D(N42), .E(n1755), .CK(clk), .Q(data_out[5]) );
  EDFFX2 \data_out_reg[4]  ( .D(N43), .E(n1755), .CK(clk), .Q(data_out[4]) );
  EDFFX2 \data_out_reg[3]  ( .D(N44), .E(n1755), .CK(clk), .Q(data_out[3]) );
  EDFFX2 \data_out_reg[2]  ( .D(N45), .E(n1755), .CK(clk), .Q(data_out[2]) );
  EDFFX2 \data_out_reg[1]  ( .D(N46), .E(n1755), .CK(clk), .Q(data_out[1]) );
  EDFFX2 \data_out_reg[0]  ( .D(N47), .E(n1755), .CK(clk), .Q(data_out[0]) );
  NOR4BX1 U2 ( .AN(wr_en), .B(index[5]), .C(index[7]), .D(index[6]), .Y(n2838)
         );
  NOR3BX2 U3 ( .AN(n2838), .B(n1408), .C(N14), .Y(n2846) );
  NOR3BX2 U4 ( .AN(n2838), .B(N14), .C(n1761), .Y(n2837) );
  NAND2X1 U5 ( .A(n2847), .B(n2846), .Y(n1) );
  NAND2X1 U6 ( .A(n2845), .B(n2846), .Y(n2) );
  NAND2X1 U7 ( .A(n2844), .B(n2846), .Y(n3) );
  NAND2X1 U8 ( .A(n2843), .B(n2846), .Y(n4) );
  NAND2X1 U9 ( .A(n2842), .B(n2846), .Y(n5) );
  NAND2X1 U10 ( .A(n2841), .B(n2846), .Y(n6) );
  NAND2X1 U11 ( .A(n2840), .B(n2846), .Y(n7) );
  NAND2X1 U12 ( .A(n2839), .B(n2846), .Y(n8) );
  NAND2X1 U13 ( .A(n2837), .B(n2847), .Y(n9) );
  NAND2X1 U14 ( .A(n2837), .B(n2845), .Y(n10) );
  NAND2X1 U15 ( .A(n2837), .B(n2844), .Y(n11) );
  NAND2X1 U16 ( .A(n2837), .B(n2843), .Y(n12) );
  NAND2X1 U17 ( .A(n2837), .B(n2842), .Y(n13) );
  NAND2X1 U18 ( .A(n2837), .B(n2841), .Y(n14) );
  NAND2X1 U19 ( .A(n2837), .B(n2840), .Y(n15) );
  NAND2X1 U20 ( .A(n2837), .B(n2839), .Y(n16) );
  NOR2X4 U21 ( .A(wr_en), .B(rst), .Y(N81) );
  CLKINVX1 U38 ( .A(n1757), .Y(n1756) );
  CLKINVX1 U39 ( .A(n1759), .Y(n1758) );
  CLKINVX1 U40 ( .A(N11), .Y(n1759) );
  CLKINVX1 U41 ( .A(N10), .Y(n1757) );
  CLKINVX1 U42 ( .A(N13), .Y(n1761) );
  CLKINVX1 U43 ( .A(rst), .Y(n1794) );
  CLKINVX1 U44 ( .A(data_in[0]), .Y(n1793) );
  CLKINVX1 U45 ( .A(data_in[1]), .Y(n1792) );
  CLKINVX1 U46 ( .A(data_in[2]), .Y(n1791) );
  CLKINVX1 U47 ( .A(data_in[3]), .Y(n1790) );
  CLKINVX1 U48 ( .A(data_in[4]), .Y(n1789) );
  CLKINVX1 U49 ( .A(data_in[5]), .Y(n1788) );
  CLKINVX1 U50 ( .A(data_in[6]), .Y(n1787) );
  CLKINVX1 U51 ( .A(data_in[7]), .Y(n1786) );
  CLKINVX1 U52 ( .A(data_in[8]), .Y(n1785) );
  CLKINVX1 U53 ( .A(data_in[9]), .Y(n1784) );
  CLKINVX1 U54 ( .A(data_in[10]), .Y(n1783) );
  CLKINVX1 U55 ( .A(data_in[11]), .Y(n1782) );
  CLKINVX1 U56 ( .A(data_in[12]), .Y(n1781) );
  CLKINVX1 U57 ( .A(data_in[13]), .Y(n1780) );
  CLKINVX1 U58 ( .A(data_in[14]), .Y(n1779) );
  CLKINVX1 U59 ( .A(data_in[15]), .Y(n1778) );
  CLKINVX1 U60 ( .A(data_in[16]), .Y(n1777) );
  CLKINVX1 U61 ( .A(data_in[17]), .Y(n1776) );
  CLKINVX1 U62 ( .A(data_in[18]), .Y(n1775) );
  CLKINVX1 U63 ( .A(data_in[19]), .Y(n1774) );
  CLKINVX1 U64 ( .A(data_in[20]), .Y(n1773) );
  CLKINVX1 U65 ( .A(data_in[21]), .Y(n1772) );
  CLKINVX1 U66 ( .A(data_in[22]), .Y(n1771) );
  CLKINVX1 U67 ( .A(data_in[23]), .Y(n1770) );
  CLKINVX1 U68 ( .A(data_in[24]), .Y(n1769) );
  CLKINVX1 U69 ( .A(data_in[25]), .Y(n1768) );
  CLKINVX1 U70 ( .A(data_in[26]), .Y(n1767) );
  CLKINVX1 U71 ( .A(data_in[27]), .Y(n1766) );
  CLKINVX1 U72 ( .A(data_in[28]), .Y(n1765) );
  CLKINVX1 U73 ( .A(data_in[29]), .Y(n1764) );
  CLKINVX1 U74 ( .A(data_in[30]), .Y(n1763) );
  CLKINVX1 U75 ( .A(data_in[31]), .Y(n1762) );
  CLKBUFX3 U76 ( .A(n1437), .Y(n1440) );
  CLKBUFX3 U77 ( .A(n1437), .Y(n1441) );
  CLKBUFX3 U78 ( .A(n1436), .Y(n1442) );
  CLKBUFX3 U79 ( .A(n1436), .Y(n1443) );
  CLKBUFX3 U80 ( .A(n1434), .Y(n1444) );
  CLKBUFX3 U81 ( .A(n1435), .Y(n1445) );
  CLKBUFX3 U82 ( .A(n1435), .Y(n1446) );
  CLKBUFX3 U83 ( .A(n1434), .Y(n1447) );
  CLKBUFX3 U84 ( .A(n1435), .Y(n1448) );
  CLKBUFX3 U85 ( .A(n1435), .Y(n1449) );
  CLKBUFX3 U86 ( .A(n1437), .Y(n1450) );
  CLKBUFX3 U87 ( .A(n1436), .Y(n1451) );
  CLKBUFX3 U88 ( .A(n1436), .Y(n1452) );
  CLKBUFX3 U89 ( .A(n1434), .Y(n1453) );
  CLKBUFX3 U90 ( .A(n1417), .Y(n1419) );
  CLKBUFX3 U91 ( .A(n1417), .Y(n1420) );
  CLKBUFX3 U92 ( .A(n1416), .Y(n1421) );
  CLKBUFX3 U93 ( .A(n1415), .Y(n1422) );
  CLKBUFX3 U94 ( .A(n1758), .Y(n1423) );
  CLKBUFX3 U95 ( .A(n1415), .Y(n1424) );
  CLKBUFX3 U96 ( .A(n1415), .Y(n1425) );
  CLKBUFX3 U97 ( .A(n1423), .Y(n1426) );
  CLKBUFX3 U98 ( .A(n1415), .Y(n1427) );
  CLKBUFX3 U99 ( .A(n1423), .Y(n1428) );
  CLKBUFX3 U100 ( .A(n1415), .Y(n1429) );
  CLKBUFX3 U101 ( .A(n1423), .Y(n1430) );
  CLKBUFX3 U102 ( .A(n1417), .Y(n1431) );
  CLKBUFX3 U103 ( .A(n1416), .Y(n1432) );
  CLKBUFX3 U104 ( .A(n1416), .Y(n1433) );
  CLKBUFX3 U105 ( .A(n1437), .Y(n1439) );
  CLKBUFX3 U106 ( .A(n1434), .Y(n1438) );
  CLKBUFX3 U107 ( .A(n1417), .Y(n1418) );
  CLKBUFX3 U108 ( .A(n1434), .Y(n1437) );
  CLKBUFX3 U109 ( .A(n1415), .Y(n1417) );
  CLKBUFX3 U110 ( .A(n1434), .Y(n1436) );
  CLKBUFX3 U111 ( .A(n1415), .Y(n1416) );
  CLKBUFX3 U112 ( .A(n1434), .Y(n1435) );
  CLKBUFX3 U113 ( .A(n1756), .Y(n1434) );
  CLKBUFX3 U114 ( .A(n1758), .Y(n1415) );
  CLKBUFX3 U115 ( .A(N13), .Y(n1408) );
  CLKBUFX3 U116 ( .A(N13), .Y(n1409) );
  CLKBUFX3 U117 ( .A(N13), .Y(n1410) );
  CLKBUFX3 U118 ( .A(N13), .Y(n1411) );
  CLKBUFX3 U119 ( .A(n1412), .Y(n1413) );
  CLKBUFX3 U120 ( .A(n1760), .Y(n1414) );
  CLKBUFX3 U121 ( .A(n1760), .Y(n1412) );
  CLKBUFX3 U122 ( .A(n1647), .Y(n1522) );
  CLKBUFX3 U123 ( .A(n1647), .Y(n1523) );
  CLKBUFX3 U124 ( .A(n1646), .Y(n1524) );
  CLKBUFX3 U125 ( .A(n1646), .Y(n1525) );
  CLKBUFX3 U126 ( .A(n1645), .Y(n1526) );
  CLKBUFX3 U127 ( .A(n1645), .Y(n1527) );
  CLKBUFX3 U128 ( .A(n1644), .Y(n1528) );
  CLKBUFX3 U129 ( .A(n1644), .Y(n1529) );
  CLKBUFX3 U130 ( .A(n1643), .Y(n1530) );
  CLKBUFX3 U131 ( .A(n1643), .Y(n1531) );
  CLKBUFX3 U132 ( .A(n1642), .Y(n1532) );
  CLKBUFX3 U133 ( .A(n1642), .Y(n1533) );
  CLKBUFX3 U134 ( .A(n1641), .Y(n1534) );
  CLKBUFX3 U135 ( .A(n1641), .Y(n1535) );
  CLKBUFX3 U136 ( .A(n1640), .Y(n1536) );
  CLKBUFX3 U137 ( .A(n1640), .Y(n1537) );
  CLKBUFX3 U138 ( .A(n1639), .Y(n1538) );
  CLKBUFX3 U139 ( .A(n1639), .Y(n1539) );
  CLKBUFX3 U140 ( .A(n1638), .Y(n1540) );
  CLKBUFX3 U141 ( .A(n1638), .Y(n1541) );
  CLKBUFX3 U142 ( .A(n1637), .Y(n1542) );
  CLKBUFX3 U143 ( .A(n1637), .Y(n1543) );
  CLKBUFX3 U144 ( .A(n1636), .Y(n1544) );
  CLKBUFX3 U145 ( .A(n1636), .Y(n1545) );
  CLKBUFX3 U146 ( .A(n1635), .Y(n1546) );
  CLKBUFX3 U147 ( .A(n1635), .Y(n1547) );
  CLKBUFX3 U148 ( .A(n1634), .Y(n1548) );
  CLKBUFX3 U149 ( .A(n1634), .Y(n1549) );
  CLKBUFX3 U150 ( .A(n1633), .Y(n1550) );
  CLKBUFX3 U151 ( .A(n1633), .Y(n1551) );
  CLKBUFX3 U152 ( .A(n1632), .Y(n1552) );
  CLKBUFX3 U153 ( .A(n1632), .Y(n1553) );
  CLKBUFX3 U154 ( .A(n1631), .Y(n1554) );
  CLKBUFX3 U155 ( .A(n1631), .Y(n1555) );
  CLKBUFX3 U156 ( .A(n1630), .Y(n1556) );
  CLKBUFX3 U157 ( .A(n1630), .Y(n1557) );
  CLKBUFX3 U158 ( .A(n1629), .Y(n1558) );
  CLKBUFX3 U159 ( .A(n1629), .Y(n1559) );
  CLKBUFX3 U160 ( .A(n1628), .Y(n1560) );
  CLKBUFX3 U161 ( .A(n1628), .Y(n1561) );
  CLKBUFX3 U162 ( .A(n1627), .Y(n1562) );
  CLKBUFX3 U163 ( .A(n1627), .Y(n1563) );
  CLKBUFX3 U164 ( .A(n1626), .Y(n1564) );
  CLKBUFX3 U165 ( .A(n1626), .Y(n1565) );
  CLKBUFX3 U166 ( .A(n1625), .Y(n1566) );
  CLKBUFX3 U167 ( .A(n1625), .Y(n1567) );
  CLKBUFX3 U168 ( .A(n1624), .Y(n1568) );
  CLKBUFX3 U169 ( .A(n1624), .Y(n1569) );
  CLKBUFX3 U170 ( .A(n1623), .Y(n1570) );
  CLKBUFX3 U171 ( .A(n1623), .Y(n1571) );
  CLKBUFX3 U172 ( .A(n1622), .Y(n1572) );
  CLKBUFX3 U173 ( .A(n1622), .Y(n1573) );
  CLKBUFX3 U174 ( .A(n1621), .Y(n1574) );
  CLKBUFX3 U175 ( .A(n1621), .Y(n1575) );
  CLKBUFX3 U176 ( .A(n1620), .Y(n1576) );
  CLKBUFX3 U177 ( .A(n1620), .Y(n1577) );
  CLKBUFX3 U178 ( .A(n1619), .Y(n1578) );
  CLKBUFX3 U179 ( .A(n1619), .Y(n1579) );
  CLKBUFX3 U180 ( .A(n1618), .Y(n1580) );
  CLKBUFX3 U181 ( .A(n1618), .Y(n1581) );
  CLKBUFX3 U182 ( .A(n1617), .Y(n1582) );
  CLKBUFX3 U183 ( .A(n1617), .Y(n1583) );
  CLKBUFX3 U184 ( .A(n1616), .Y(n1584) );
  CLKBUFX3 U185 ( .A(n1616), .Y(n1585) );
  CLKBUFX3 U186 ( .A(n1615), .Y(n1586) );
  CLKBUFX3 U187 ( .A(n1615), .Y(n1587) );
  CLKBUFX3 U188 ( .A(n1614), .Y(n1588) );
  CLKBUFX3 U189 ( .A(n1614), .Y(n1589) );
  CLKBUFX3 U190 ( .A(n1613), .Y(n1590) );
  CLKBUFX3 U191 ( .A(n1613), .Y(n1591) );
  CLKBUFX3 U192 ( .A(n1612), .Y(n1592) );
  CLKBUFX3 U193 ( .A(n1612), .Y(n1593) );
  CLKBUFX3 U194 ( .A(n1611), .Y(n1594) );
  CLKBUFX3 U195 ( .A(n1611), .Y(n1595) );
  CLKBUFX3 U196 ( .A(n1610), .Y(n1596) );
  CLKBUFX3 U197 ( .A(n1610), .Y(n1597) );
  CLKBUFX3 U198 ( .A(n1609), .Y(n1598) );
  CLKBUFX3 U199 ( .A(n1609), .Y(n1599) );
  CLKBUFX3 U200 ( .A(n1608), .Y(n1600) );
  CLKBUFX3 U201 ( .A(n1608), .Y(n1601) );
  CLKBUFX3 U202 ( .A(n1658), .Y(n1602) );
  CLKBUFX3 U203 ( .A(n1646), .Y(n1603) );
  CLKBUFX3 U204 ( .A(n1658), .Y(n1604) );
  CLKBUFX3 U205 ( .A(n1647), .Y(n1605) );
  CLKBUFX3 U206 ( .A(n1658), .Y(n1606) );
  CLKBUFX3 U207 ( .A(n1), .Y(n1754) );
  CLKBUFX3 U208 ( .A(n1), .Y(n1753) );
  CLKBUFX3 U209 ( .A(n2), .Y(n1750) );
  CLKBUFX3 U210 ( .A(n3), .Y(n1747) );
  CLKBUFX3 U211 ( .A(n4), .Y(n1744) );
  CLKBUFX3 U212 ( .A(n6), .Y(n1738) );
  CLKBUFX3 U213 ( .A(n7), .Y(n1735) );
  CLKBUFX3 U214 ( .A(n8), .Y(n1732) );
  CLKBUFX3 U215 ( .A(n9), .Y(n1729) );
  CLKBUFX3 U216 ( .A(n10), .Y(n1726) );
  CLKBUFX3 U217 ( .A(n11), .Y(n1723) );
  CLKBUFX3 U218 ( .A(n12), .Y(n1720) );
  CLKBUFX3 U219 ( .A(n14), .Y(n1714) );
  CLKBUFX3 U220 ( .A(n15), .Y(n1711) );
  CLKBUFX3 U221 ( .A(n16), .Y(n1708) );
  CLKBUFX3 U222 ( .A(n2836), .Y(n1705) );
  CLKBUFX3 U223 ( .A(n2834), .Y(n1702) );
  CLKBUFX3 U224 ( .A(n2833), .Y(n1699) );
  CLKBUFX3 U225 ( .A(n2832), .Y(n1696) );
  CLKBUFX3 U226 ( .A(n2831), .Y(n1693) );
  CLKBUFX3 U227 ( .A(n2830), .Y(n1690) );
  CLKBUFX3 U228 ( .A(n2829), .Y(n1687) );
  CLKBUFX3 U229 ( .A(n2828), .Y(n1684) );
  CLKBUFX3 U230 ( .A(n2827), .Y(n1681) );
  CLKBUFX3 U231 ( .A(n2825), .Y(n1678) );
  CLKBUFX3 U232 ( .A(n2824), .Y(n1675) );
  CLKBUFX3 U233 ( .A(n2823), .Y(n1672) );
  CLKBUFX3 U234 ( .A(n2822), .Y(n1669) );
  CLKBUFX3 U235 ( .A(n2821), .Y(n1666) );
  CLKBUFX3 U236 ( .A(n2820), .Y(n1663) );
  CLKBUFX3 U237 ( .A(n2819), .Y(n1660) );
  CLKBUFX3 U238 ( .A(n1), .Y(n1752) );
  CLKBUFX3 U239 ( .A(n2), .Y(n1751) );
  CLKBUFX3 U240 ( .A(n3), .Y(n1748) );
  CLKBUFX3 U241 ( .A(n4), .Y(n1745) );
  CLKBUFX3 U242 ( .A(n5), .Y(n1742) );
  CLKBUFX3 U243 ( .A(n6), .Y(n1739) );
  CLKBUFX3 U244 ( .A(n7), .Y(n1736) );
  CLKBUFX3 U245 ( .A(n8), .Y(n1733) );
  CLKBUFX3 U246 ( .A(n9), .Y(n1730) );
  CLKBUFX3 U247 ( .A(n10), .Y(n1727) );
  CLKBUFX3 U248 ( .A(n11), .Y(n1724) );
  CLKBUFX3 U249 ( .A(n12), .Y(n1721) );
  CLKBUFX3 U250 ( .A(n13), .Y(n1718) );
  CLKBUFX3 U251 ( .A(n14), .Y(n1715) );
  CLKBUFX3 U252 ( .A(n15), .Y(n1712) );
  CLKBUFX3 U253 ( .A(n16), .Y(n1709) );
  CLKBUFX3 U254 ( .A(n2836), .Y(n1706) );
  CLKBUFX3 U255 ( .A(n2834), .Y(n1703) );
  CLKBUFX3 U256 ( .A(n2833), .Y(n1700) );
  CLKBUFX3 U257 ( .A(n2832), .Y(n1697) );
  CLKBUFX3 U258 ( .A(n2831), .Y(n1694) );
  CLKBUFX3 U259 ( .A(n2830), .Y(n1691) );
  CLKBUFX3 U260 ( .A(n2829), .Y(n1688) );
  CLKBUFX3 U261 ( .A(n2828), .Y(n1685) );
  CLKBUFX3 U262 ( .A(n2827), .Y(n1682) );
  CLKBUFX3 U263 ( .A(n2825), .Y(n1679) );
  CLKBUFX3 U264 ( .A(n2824), .Y(n1676) );
  CLKBUFX3 U265 ( .A(n2823), .Y(n1673) );
  CLKBUFX3 U266 ( .A(n2822), .Y(n1670) );
  CLKBUFX3 U267 ( .A(n2821), .Y(n1667) );
  CLKBUFX3 U268 ( .A(n2820), .Y(n1664) );
  CLKBUFX3 U269 ( .A(n2819), .Y(n1661) );
  CLKBUFX3 U270 ( .A(n2), .Y(n1749) );
  CLKBUFX3 U271 ( .A(n3), .Y(n1746) );
  CLKBUFX3 U272 ( .A(n4), .Y(n1743) );
  CLKBUFX3 U273 ( .A(n5), .Y(n1740) );
  CLKBUFX3 U274 ( .A(n5), .Y(n1741) );
  CLKBUFX3 U275 ( .A(n6), .Y(n1737) );
  CLKBUFX3 U276 ( .A(n7), .Y(n1734) );
  CLKBUFX3 U277 ( .A(n8), .Y(n1731) );
  CLKBUFX3 U278 ( .A(n9), .Y(n1728) );
  CLKBUFX3 U279 ( .A(n10), .Y(n1725) );
  CLKBUFX3 U280 ( .A(n11), .Y(n1722) );
  CLKBUFX3 U281 ( .A(n12), .Y(n1719) );
  CLKBUFX3 U282 ( .A(n13), .Y(n1716) );
  CLKBUFX3 U283 ( .A(n13), .Y(n1717) );
  CLKBUFX3 U284 ( .A(n14), .Y(n1713) );
  CLKBUFX3 U285 ( .A(n15), .Y(n1710) );
  CLKBUFX3 U286 ( .A(n16), .Y(n1707) );
  CLKBUFX3 U287 ( .A(n2836), .Y(n1704) );
  CLKBUFX3 U288 ( .A(n2834), .Y(n1701) );
  CLKBUFX3 U289 ( .A(n2833), .Y(n1698) );
  CLKBUFX3 U290 ( .A(n2832), .Y(n1695) );
  CLKBUFX3 U291 ( .A(n2831), .Y(n1692) );
  CLKBUFX3 U292 ( .A(n2830), .Y(n1689) );
  CLKBUFX3 U293 ( .A(n2829), .Y(n1686) );
  CLKBUFX3 U294 ( .A(n2828), .Y(n1683) );
  CLKBUFX3 U295 ( .A(n2827), .Y(n1680) );
  CLKBUFX3 U296 ( .A(n2825), .Y(n1677) );
  CLKBUFX3 U297 ( .A(n2824), .Y(n1674) );
  CLKBUFX3 U298 ( .A(n2823), .Y(n1671) );
  CLKBUFX3 U299 ( .A(n2822), .Y(n1668) );
  CLKBUFX3 U300 ( .A(n2821), .Y(n1665) );
  CLKBUFX3 U301 ( .A(n2820), .Y(n1662) );
  CLKBUFX3 U302 ( .A(n2819), .Y(n1659) );
  CLKBUFX3 U303 ( .A(n1521), .Y(n1607) );
  CLKBUFX3 U304 ( .A(N14), .Y(n1406) );
  CLKBUFX3 U305 ( .A(N14), .Y(n1407) );
  NOR3X1 U306 ( .A(n1758), .B(n1760), .C(n1756), .Y(n2847) );
  NOR3X1 U307 ( .A(n1758), .B(n1760), .C(n1757), .Y(n2845) );
  NOR3X1 U308 ( .A(n1756), .B(n1760), .C(n1759), .Y(n2844) );
  NOR3X1 U309 ( .A(n1757), .B(n1760), .C(n1759), .Y(n2843) );
  AND3X2 U310 ( .A(n1760), .B(n1757), .C(n1759), .Y(n2842) );
  AND3X2 U311 ( .A(n1760), .B(n1756), .C(n1759), .Y(n2841) );
  AND3X2 U312 ( .A(n1760), .B(n1758), .C(n1757), .Y(n2840) );
  AND3X2 U313 ( .A(n1760), .B(n1758), .C(n1756), .Y(n2839) );
  CLKBUFX3 U314 ( .A(n1648), .Y(n1647) );
  CLKBUFX3 U315 ( .A(n1648), .Y(n1646) );
  CLKBUFX3 U316 ( .A(n1648), .Y(n1645) );
  CLKBUFX3 U317 ( .A(n1648), .Y(n1644) );
  CLKBUFX3 U318 ( .A(n1649), .Y(n1643) );
  CLKBUFX3 U319 ( .A(n1649), .Y(n1642) );
  CLKBUFX3 U320 ( .A(n1649), .Y(n1641) );
  CLKBUFX3 U321 ( .A(n1649), .Y(n1640) );
  CLKBUFX3 U322 ( .A(n1650), .Y(n1639) );
  CLKBUFX3 U323 ( .A(n1650), .Y(n1638) );
  CLKBUFX3 U324 ( .A(n1650), .Y(n1637) );
  CLKBUFX3 U325 ( .A(n1650), .Y(n1636) );
  CLKBUFX3 U326 ( .A(n1651), .Y(n1635) );
  CLKBUFX3 U327 ( .A(n1651), .Y(n1634) );
  CLKBUFX3 U328 ( .A(n1651), .Y(n1633) );
  CLKBUFX3 U329 ( .A(n1651), .Y(n1632) );
  CLKBUFX3 U330 ( .A(n1652), .Y(n1631) );
  CLKBUFX3 U331 ( .A(n1652), .Y(n1630) );
  CLKBUFX3 U332 ( .A(n1652), .Y(n1629) );
  CLKBUFX3 U333 ( .A(n1652), .Y(n1628) );
  CLKBUFX3 U334 ( .A(n1653), .Y(n1627) );
  CLKBUFX3 U335 ( .A(n1653), .Y(n1626) );
  CLKBUFX3 U336 ( .A(n1653), .Y(n1625) );
  CLKBUFX3 U337 ( .A(n1653), .Y(n1624) );
  CLKBUFX3 U338 ( .A(n1654), .Y(n1623) );
  CLKBUFX3 U339 ( .A(n1654), .Y(n1622) );
  CLKBUFX3 U340 ( .A(n1654), .Y(n1621) );
  CLKBUFX3 U341 ( .A(n1654), .Y(n1620) );
  CLKBUFX3 U342 ( .A(n1655), .Y(n1619) );
  CLKBUFX3 U343 ( .A(n1655), .Y(n1618) );
  CLKBUFX3 U344 ( .A(n1655), .Y(n1617) );
  CLKBUFX3 U345 ( .A(n1655), .Y(n1616) );
  CLKBUFX3 U346 ( .A(n1656), .Y(n1615) );
  CLKBUFX3 U347 ( .A(n1656), .Y(n1614) );
  CLKBUFX3 U348 ( .A(n1656), .Y(n1613) );
  CLKBUFX3 U349 ( .A(n1656), .Y(n1612) );
  CLKBUFX3 U350 ( .A(n1657), .Y(n1611) );
  CLKBUFX3 U351 ( .A(n1657), .Y(n1610) );
  CLKBUFX3 U352 ( .A(n1657), .Y(n1609) );
  CLKBUFX3 U353 ( .A(n1657), .Y(n1608) );
  CLKBUFX3 U354 ( .A(N12), .Y(n1760) );
  NAND2X1 U355 ( .A(n2835), .B(n2847), .Y(n2836) );
  NAND2X1 U356 ( .A(n2835), .B(n2845), .Y(n2834) );
  NAND2X1 U357 ( .A(n2835), .B(n2844), .Y(n2833) );
  NAND2X1 U358 ( .A(n2835), .B(n2843), .Y(n2832) );
  NAND2X1 U359 ( .A(n2826), .B(n2847), .Y(n2827) );
  NAND2X1 U360 ( .A(n2826), .B(n2845), .Y(n2825) );
  NAND2X1 U361 ( .A(n2826), .B(n2844), .Y(n2824) );
  NAND2X1 U362 ( .A(n2826), .B(n2843), .Y(n2823) );
  NAND2X1 U363 ( .A(n2835), .B(n2842), .Y(n2831) );
  NAND2X1 U364 ( .A(n2835), .B(n2841), .Y(n2830) );
  NAND2X1 U365 ( .A(n2835), .B(n2840), .Y(n2829) );
  NAND2X1 U366 ( .A(n2835), .B(n2839), .Y(n2828) );
  NAND2X1 U367 ( .A(n2826), .B(n2842), .Y(n2822) );
  NAND2X1 U368 ( .A(n2826), .B(n2841), .Y(n2821) );
  NAND2X1 U369 ( .A(n2826), .B(n2840), .Y(n2820) );
  NAND2X1 U370 ( .A(n2826), .B(n2839), .Y(n2819) );
  CLKBUFX3 U371 ( .A(n1518), .Y(n1648) );
  CLKBUFX3 U372 ( .A(n1518), .Y(n1649) );
  CLKBUFX3 U373 ( .A(n1518), .Y(n1650) );
  CLKBUFX3 U374 ( .A(n1519), .Y(n1651) );
  CLKBUFX3 U375 ( .A(n1519), .Y(n1652) );
  CLKBUFX3 U376 ( .A(n1519), .Y(n1653) );
  CLKBUFX3 U377 ( .A(n1520), .Y(n1654) );
  CLKBUFX3 U378 ( .A(n1520), .Y(n1655) );
  CLKBUFX3 U379 ( .A(n1520), .Y(n1656) );
  CLKBUFX3 U380 ( .A(n1521), .Y(n1657) );
  CLKBUFX3 U381 ( .A(n1521), .Y(n1658) );
  CLKBUFX3 U382 ( .A(N81), .Y(n1755) );
  AND3X2 U383 ( .A(n2838), .B(n1761), .C(N14), .Y(n2835) );
  AND3X2 U384 ( .A(n1411), .B(n2838), .C(N14), .Y(n2826) );
  CLKBUFX3 U385 ( .A(n1794), .Y(n1518) );
  CLKBUFX3 U386 ( .A(n1794), .Y(n1519) );
  CLKBUFX3 U387 ( .A(n1794), .Y(n1520) );
  CLKBUFX3 U388 ( .A(n1794), .Y(n1521) );
  CLKBUFX3 U389 ( .A(n1793), .Y(n1517) );
  CLKBUFX3 U390 ( .A(n1792), .Y(n1515) );
  CLKBUFX3 U391 ( .A(n1791), .Y(n1513) );
  CLKBUFX3 U392 ( .A(n1790), .Y(n1511) );
  CLKBUFX3 U393 ( .A(n1789), .Y(n1509) );
  CLKBUFX3 U394 ( .A(n1788), .Y(n1507) );
  CLKBUFX3 U395 ( .A(n1787), .Y(n1505) );
  CLKBUFX3 U396 ( .A(n1786), .Y(n1503) );
  CLKBUFX3 U397 ( .A(n1785), .Y(n1501) );
  CLKBUFX3 U398 ( .A(n1784), .Y(n1499) );
  CLKBUFX3 U399 ( .A(n1783), .Y(n1497) );
  CLKBUFX3 U400 ( .A(n1782), .Y(n1495) );
  CLKBUFX3 U401 ( .A(n1781), .Y(n1493) );
  CLKBUFX3 U402 ( .A(n1780), .Y(n1491) );
  CLKBUFX3 U403 ( .A(n1779), .Y(n1489) );
  CLKBUFX3 U404 ( .A(n1778), .Y(n1487) );
  CLKBUFX3 U405 ( .A(n1777), .Y(n1485) );
  CLKBUFX3 U406 ( .A(n1776), .Y(n1483) );
  CLKBUFX3 U407 ( .A(n1775), .Y(n1481) );
  CLKBUFX3 U408 ( .A(n1774), .Y(n1479) );
  CLKBUFX3 U409 ( .A(n1773), .Y(n1477) );
  CLKBUFX3 U410 ( .A(n1772), .Y(n1475) );
  CLKBUFX3 U411 ( .A(n1771), .Y(n1473) );
  CLKBUFX3 U412 ( .A(n1770), .Y(n1471) );
  CLKBUFX3 U413 ( .A(n1769), .Y(n1469) );
  CLKBUFX3 U414 ( .A(n1768), .Y(n1467) );
  CLKBUFX3 U415 ( .A(n1767), .Y(n1465) );
  CLKBUFX3 U416 ( .A(n1766), .Y(n1463) );
  CLKBUFX3 U417 ( .A(n1765), .Y(n1461) );
  CLKBUFX3 U418 ( .A(n1764), .Y(n1459) );
  CLKBUFX3 U419 ( .A(n1763), .Y(n1457) );
  CLKBUFX3 U420 ( .A(n1762), .Y(n1455) );
  CLKBUFX3 U421 ( .A(n1793), .Y(n1516) );
  CLKBUFX3 U422 ( .A(n1792), .Y(n1514) );
  CLKBUFX3 U423 ( .A(n1791), .Y(n1512) );
  CLKBUFX3 U424 ( .A(n1790), .Y(n1510) );
  CLKBUFX3 U425 ( .A(n1789), .Y(n1508) );
  CLKBUFX3 U426 ( .A(n1788), .Y(n1506) );
  CLKBUFX3 U427 ( .A(n1787), .Y(n1504) );
  CLKBUFX3 U428 ( .A(n1786), .Y(n1502) );
  CLKBUFX3 U429 ( .A(n1785), .Y(n1500) );
  CLKBUFX3 U430 ( .A(n1784), .Y(n1498) );
  CLKBUFX3 U431 ( .A(n1783), .Y(n1496) );
  CLKBUFX3 U432 ( .A(n1782), .Y(n1494) );
  CLKBUFX3 U433 ( .A(n1781), .Y(n1492) );
  CLKBUFX3 U434 ( .A(n1780), .Y(n1490) );
  CLKBUFX3 U435 ( .A(n1779), .Y(n1488) );
  CLKBUFX3 U436 ( .A(n1778), .Y(n1486) );
  CLKBUFX3 U437 ( .A(n1777), .Y(n1484) );
  CLKBUFX3 U438 ( .A(n1776), .Y(n1482) );
  CLKBUFX3 U439 ( .A(n1775), .Y(n1480) );
  CLKBUFX3 U440 ( .A(n1774), .Y(n1478) );
  CLKBUFX3 U441 ( .A(n1773), .Y(n1476) );
  CLKBUFX3 U442 ( .A(n1772), .Y(n1474) );
  CLKBUFX3 U443 ( .A(n1771), .Y(n1472) );
  CLKBUFX3 U444 ( .A(n1770), .Y(n1470) );
  CLKBUFX3 U445 ( .A(n1769), .Y(n1468) );
  CLKBUFX3 U446 ( .A(n1768), .Y(n1466) );
  CLKBUFX3 U447 ( .A(n1767), .Y(n1464) );
  CLKBUFX3 U448 ( .A(n1766), .Y(n1462) );
  CLKBUFX3 U449 ( .A(n1765), .Y(n1460) );
  CLKBUFX3 U450 ( .A(n1764), .Y(n1458) );
  CLKBUFX3 U451 ( .A(n1763), .Y(n1456) );
  CLKBUFX3 U452 ( .A(n1762), .Y(n1454) );
  MX4X1 U453 ( .A(\gbuff[4][0] ), .B(\gbuff[5][0] ), .C(\gbuff[6][0] ), .D(
        \gbuff[7][0] ), .S0(n1438), .S1(n1424), .Y(n39) );
  MX4X1 U454 ( .A(\gbuff[20][0] ), .B(\gbuff[21][0] ), .C(\gbuff[22][0] ), .D(
        \gbuff[23][0] ), .S0(n1438), .S1(n1425), .Y(n35) );
  MX4X1 U455 ( .A(\gbuff[4][1] ), .B(\gbuff[5][1] ), .C(\gbuff[6][1] ), .D(
        \gbuff[7][1] ), .S0(n1439), .S1(n1418), .Y(n49) );
  MX4X1 U456 ( .A(\gbuff[20][1] ), .B(\gbuff[21][1] ), .C(\gbuff[22][1] ), .D(
        \gbuff[23][1] ), .S0(n1439), .S1(n1418), .Y(n45) );
  MX4X1 U457 ( .A(\gbuff[4][2] ), .B(\gbuff[5][2] ), .C(\gbuff[6][2] ), .D(
        \gbuff[7][2] ), .S0(n1440), .S1(n1419), .Y(n59) );
  MX4X1 U458 ( .A(\gbuff[20][2] ), .B(\gbuff[21][2] ), .C(\gbuff[22][2] ), .D(
        \gbuff[23][2] ), .S0(n1439), .S1(n1418), .Y(n55) );
  MX4X1 U459 ( .A(\gbuff[4][3] ), .B(\gbuff[5][3] ), .C(\gbuff[6][3] ), .D(
        \gbuff[7][3] ), .S0(n1440), .S1(n1419), .Y(n69) );
  MX4X1 U460 ( .A(\gbuff[20][3] ), .B(\gbuff[21][3] ), .C(\gbuff[22][3] ), .D(
        \gbuff[23][3] ), .S0(n1440), .S1(n1419), .Y(n65) );
  MX4X1 U461 ( .A(\gbuff[4][4] ), .B(\gbuff[5][4] ), .C(\gbuff[6][4] ), .D(
        \gbuff[7][4] ), .S0(n1441), .S1(n1420), .Y(n79) );
  MX4X1 U462 ( .A(\gbuff[20][4] ), .B(\gbuff[21][4] ), .C(\gbuff[22][4] ), .D(
        \gbuff[23][4] ), .S0(n1440), .S1(n1419), .Y(n75) );
  MX4X1 U463 ( .A(\gbuff[4][5] ), .B(\gbuff[5][5] ), .C(\gbuff[6][5] ), .D(
        \gbuff[7][5] ), .S0(n1441), .S1(n1420), .Y(n89) );
  MX4X1 U464 ( .A(\gbuff[20][5] ), .B(\gbuff[21][5] ), .C(\gbuff[22][5] ), .D(
        \gbuff[23][5] ), .S0(n1441), .S1(n1420), .Y(n85) );
  MX4X1 U465 ( .A(\gbuff[4][6] ), .B(\gbuff[5][6] ), .C(\gbuff[6][6] ), .D(
        \gbuff[7][6] ), .S0(n1442), .S1(n1421), .Y(n99) );
  MX4X1 U466 ( .A(\gbuff[20][6] ), .B(\gbuff[21][6] ), .C(\gbuff[22][6] ), .D(
        \gbuff[23][6] ), .S0(n1442), .S1(n1421), .Y(n95) );
  MX4X1 U467 ( .A(\gbuff[4][7] ), .B(\gbuff[5][7] ), .C(\gbuff[6][7] ), .D(
        \gbuff[7][7] ), .S0(n1443), .S1(n1431), .Y(n119) );
  MX4X1 U468 ( .A(\gbuff[20][7] ), .B(\gbuff[21][7] ), .C(\gbuff[22][7] ), .D(
        \gbuff[23][7] ), .S0(n1442), .S1(n1421), .Y(n110) );
  MX4X1 U469 ( .A(\gbuff[4][8] ), .B(\gbuff[5][8] ), .C(\gbuff[6][8] ), .D(
        \gbuff[7][8] ), .S0(n1443), .S1(n1415), .Y(n1172) );
  MX4X1 U470 ( .A(\gbuff[20][8] ), .B(\gbuff[21][8] ), .C(\gbuff[22][8] ), .D(
        \gbuff[23][8] ), .S0(n1443), .S1(n1415), .Y(n126) );
  MX4X1 U471 ( .A(\gbuff[4][9] ), .B(\gbuff[5][9] ), .C(\gbuff[6][9] ), .D(
        \gbuff[7][9] ), .S0(n1444), .S1(n1422), .Y(n1182) );
  MX4X1 U472 ( .A(\gbuff[20][9] ), .B(\gbuff[21][9] ), .C(\gbuff[22][9] ), .D(
        \gbuff[23][9] ), .S0(n1444), .S1(n1422), .Y(n1178) );
  MX4X1 U473 ( .A(\gbuff[4][10] ), .B(\gbuff[5][10] ), .C(\gbuff[6][10] ), .D(
        \gbuff[7][10] ), .S0(n1444), .S1(n1422), .Y(n1192) );
  MX4X1 U474 ( .A(\gbuff[20][10] ), .B(\gbuff[21][10] ), .C(\gbuff[22][10] ), 
        .D(\gbuff[23][10] ), .S0(n1444), .S1(n1422), .Y(n1188) );
  MX4X1 U475 ( .A(\gbuff[4][11] ), .B(\gbuff[5][11] ), .C(\gbuff[6][11] ), .D(
        \gbuff[7][11] ), .S0(n1437), .S1(n1423), .Y(n1202) );
  MX4X1 U476 ( .A(\gbuff[20][11] ), .B(\gbuff[21][11] ), .C(\gbuff[22][11] ), 
        .D(\gbuff[23][11] ), .S0(n1436), .S1(n1423), .Y(n1198) );
  MX4X1 U477 ( .A(\gbuff[4][12] ), .B(\gbuff[5][12] ), .C(\gbuff[6][12] ), .D(
        \gbuff[7][12] ), .S0(n1445), .S1(n1424), .Y(n1212) );
  MX4X1 U478 ( .A(\gbuff[20][12] ), .B(\gbuff[21][12] ), .C(\gbuff[22][12] ), 
        .D(\gbuff[23][12] ), .S0(n1435), .S1(n1423), .Y(n1208) );
  MX4X1 U479 ( .A(\gbuff[4][13] ), .B(\gbuff[5][13] ), .C(\gbuff[6][13] ), .D(
        \gbuff[7][13] ), .S0(n1445), .S1(n1424), .Y(n1222) );
  MX4X1 U480 ( .A(\gbuff[20][13] ), .B(\gbuff[21][13] ), .C(\gbuff[22][13] ), 
        .D(\gbuff[23][13] ), .S0(n1445), .S1(n1424), .Y(n1218) );
  MX4X1 U481 ( .A(\gbuff[4][14] ), .B(\gbuff[5][14] ), .C(\gbuff[6][14] ), .D(
        \gbuff[7][14] ), .S0(n1446), .S1(n1425), .Y(n1232) );
  MX4X1 U482 ( .A(\gbuff[20][14] ), .B(\gbuff[21][14] ), .C(\gbuff[22][14] ), 
        .D(\gbuff[23][14] ), .S0(n1446), .S1(n1425), .Y(n1228) );
  MX4X1 U483 ( .A(\gbuff[4][15] ), .B(\gbuff[5][15] ), .C(\gbuff[6][15] ), .D(
        \gbuff[7][15] ), .S0(n1447), .S1(n1426), .Y(n1242) );
  MX4X1 U484 ( .A(\gbuff[20][15] ), .B(\gbuff[21][15] ), .C(\gbuff[22][15] ), 
        .D(\gbuff[23][15] ), .S0(n1446), .S1(n1425), .Y(n1238) );
  MX4X1 U485 ( .A(\gbuff[4][16] ), .B(\gbuff[5][16] ), .C(\gbuff[6][16] ), .D(
        \gbuff[7][16] ), .S0(n1447), .S1(n1426), .Y(n1252) );
  MX4X1 U486 ( .A(\gbuff[20][16] ), .B(\gbuff[21][16] ), .C(\gbuff[22][16] ), 
        .D(\gbuff[23][16] ), .S0(n1447), .S1(n1426), .Y(n1248) );
  MX4X1 U487 ( .A(\gbuff[4][17] ), .B(\gbuff[5][17] ), .C(\gbuff[6][17] ), .D(
        \gbuff[7][17] ), .S0(n1436), .S1(n1427), .Y(n1262) );
  MX4X1 U488 ( .A(\gbuff[20][17] ), .B(\gbuff[21][17] ), .C(\gbuff[22][17] ), 
        .D(\gbuff[23][17] ), .S0(n1447), .S1(n1426), .Y(n1258) );
  MX4X1 U489 ( .A(\gbuff[4][18] ), .B(\gbuff[5][18] ), .C(\gbuff[6][18] ), .D(
        \gbuff[7][18] ), .S0(n1435), .S1(n1427), .Y(n1272) );
  MX4X1 U490 ( .A(\gbuff[20][18] ), .B(\gbuff[21][18] ), .C(\gbuff[22][18] ), 
        .D(\gbuff[23][18] ), .S0(n1437), .S1(n1427), .Y(n1268) );
  MX4X1 U491 ( .A(\gbuff[4][19] ), .B(\gbuff[5][19] ), .C(\gbuff[6][19] ), .D(
        \gbuff[7][19] ), .S0(n1436), .S1(n1428), .Y(n1282) );
  MX4X1 U492 ( .A(\gbuff[20][19] ), .B(\gbuff[21][19] ), .C(\gbuff[22][19] ), 
        .D(\gbuff[23][19] ), .S0(n1437), .S1(n1428), .Y(n1278) );
  MX4X1 U493 ( .A(\gbuff[4][20] ), .B(\gbuff[5][20] ), .C(\gbuff[6][20] ), .D(
        \gbuff[7][20] ), .S0(n1448), .S1(n1429), .Y(n1292) );
  MX4X1 U494 ( .A(\gbuff[20][20] ), .B(\gbuff[21][20] ), .C(\gbuff[22][20] ), 
        .D(\gbuff[23][20] ), .S0(n1435), .S1(n1428), .Y(n1288) );
  MX4X1 U495 ( .A(\gbuff[4][21] ), .B(\gbuff[5][21] ), .C(\gbuff[6][21] ), .D(
        \gbuff[7][21] ), .S0(n1448), .S1(n1429), .Y(n1302) );
  MX4X1 U496 ( .A(\gbuff[20][21] ), .B(\gbuff[21][21] ), .C(\gbuff[22][21] ), 
        .D(\gbuff[23][21] ), .S0(n1448), .S1(n1429), .Y(n1298) );
  MX4X1 U497 ( .A(\gbuff[4][22] ), .B(\gbuff[5][22] ), .C(\gbuff[6][22] ), .D(
        \gbuff[7][22] ), .S0(N10), .S1(n1430), .Y(n1312) );
  MX4X1 U498 ( .A(\gbuff[20][22] ), .B(\gbuff[21][22] ), .C(\gbuff[22][22] ), 
        .D(\gbuff[23][22] ), .S0(n1434), .S1(n1430), .Y(n1308) );
  MX4X1 U499 ( .A(\gbuff[4][23] ), .B(\gbuff[5][23] ), .C(\gbuff[6][23] ), .D(
        \gbuff[7][23] ), .S0(n1434), .S1(n1430), .Y(n1322) );
  MX4X1 U500 ( .A(\gbuff[20][23] ), .B(\gbuff[21][23] ), .C(\gbuff[22][23] ), 
        .D(\gbuff[23][23] ), .S0(n1434), .S1(n1430), .Y(n1318) );
  MX4X1 U501 ( .A(\gbuff[4][24] ), .B(\gbuff[5][24] ), .C(\gbuff[6][24] ), .D(
        \gbuff[7][24] ), .S0(n1449), .S1(n1428), .Y(n1332) );
  MX4X1 U502 ( .A(\gbuff[20][24] ), .B(\gbuff[21][24] ), .C(\gbuff[22][24] ), 
        .D(\gbuff[23][24] ), .S0(n1449), .S1(n1430), .Y(n1328) );
  MX4X1 U503 ( .A(\gbuff[4][25] ), .B(\gbuff[5][25] ), .C(\gbuff[6][25] ), .D(
        \gbuff[7][25] ), .S0(n1450), .S1(n1431), .Y(n1342) );
  MX4X1 U504 ( .A(\gbuff[20][25] ), .B(\gbuff[21][25] ), .C(\gbuff[22][25] ), 
        .D(\gbuff[23][25] ), .S0(n1449), .S1(n1415), .Y(n1338) );
  MX4X1 U505 ( .A(\gbuff[4][26] ), .B(\gbuff[5][26] ), .C(\gbuff[6][26] ), .D(
        \gbuff[7][26] ), .S0(n1450), .S1(n1431), .Y(n1352) );
  MX4X1 U506 ( .A(\gbuff[20][26] ), .B(\gbuff[21][26] ), .C(\gbuff[22][26] ), 
        .D(\gbuff[23][26] ), .S0(n1450), .S1(n1431), .Y(n1348) );
  MX4X1 U507 ( .A(\gbuff[4][27] ), .B(\gbuff[5][27] ), .C(\gbuff[6][27] ), .D(
        \gbuff[7][27] ), .S0(n1451), .S1(n1432), .Y(n1362) );
  MX4X1 U508 ( .A(\gbuff[20][27] ), .B(\gbuff[21][27] ), .C(\gbuff[22][27] ), 
        .D(\gbuff[23][27] ), .S0(n1451), .S1(n1432), .Y(n1358) );
  MX4X1 U509 ( .A(\gbuff[4][28] ), .B(\gbuff[5][28] ), .C(\gbuff[6][28] ), .D(
        \gbuff[7][28] ), .S0(n1452), .S1(n1433), .Y(n1372) );
  MX4X1 U510 ( .A(\gbuff[20][28] ), .B(\gbuff[21][28] ), .C(\gbuff[22][28] ), 
        .D(\gbuff[23][28] ), .S0(n1451), .S1(n1432), .Y(n1368) );
  MX4X1 U511 ( .A(\gbuff[4][29] ), .B(\gbuff[5][29] ), .C(\gbuff[6][29] ), .D(
        \gbuff[7][29] ), .S0(n1452), .S1(n1433), .Y(n1382) );
  MX4X1 U512 ( .A(\gbuff[20][29] ), .B(\gbuff[21][29] ), .C(\gbuff[22][29] ), 
        .D(\gbuff[23][29] ), .S0(n1452), .S1(n1433), .Y(n1378) );
  MX4X1 U513 ( .A(\gbuff[4][30] ), .B(\gbuff[5][30] ), .C(\gbuff[6][30] ), .D(
        \gbuff[7][30] ), .S0(n1453), .S1(n1425), .Y(n1392) );
  MX4X1 U514 ( .A(\gbuff[20][30] ), .B(\gbuff[21][30] ), .C(\gbuff[22][30] ), 
        .D(\gbuff[23][30] ), .S0(n1452), .S1(n1433), .Y(n1388) );
  MX4X1 U515 ( .A(\gbuff[4][31] ), .B(\gbuff[5][31] ), .C(\gbuff[6][31] ), .D(
        \gbuff[7][31] ), .S0(n1453), .S1(n1424), .Y(n1402) );
  MX4X1 U516 ( .A(\gbuff[20][31] ), .B(\gbuff[21][31] ), .C(\gbuff[22][31] ), 
        .D(\gbuff[23][31] ), .S0(n1453), .S1(n1422), .Y(n1398) );
  MX4X1 U517 ( .A(\gbuff[0][0] ), .B(\gbuff[1][0] ), .C(\gbuff[2][0] ), .D(
        \gbuff[3][0] ), .S0(n1438), .S1(n1422), .Y(n40) );
  MX4X1 U518 ( .A(\gbuff[16][0] ), .B(\gbuff[17][0] ), .C(\gbuff[18][0] ), .D(
        \gbuff[19][0] ), .S0(n1438), .S1(n1427), .Y(n36) );
  MX4X1 U519 ( .A(\gbuff[0][1] ), .B(\gbuff[1][1] ), .C(\gbuff[2][1] ), .D(
        \gbuff[3][1] ), .S0(n1439), .S1(n1418), .Y(n50) );
  MX4X1 U520 ( .A(\gbuff[16][1] ), .B(\gbuff[17][1] ), .C(\gbuff[18][1] ), .D(
        \gbuff[19][1] ), .S0(n1439), .S1(n1418), .Y(n46) );
  MX4X1 U521 ( .A(\gbuff[0][2] ), .B(\gbuff[1][2] ), .C(\gbuff[2][2] ), .D(
        \gbuff[3][2] ), .S0(n1440), .S1(n1419), .Y(n60) );
  MX4X1 U522 ( .A(\gbuff[16][2] ), .B(\gbuff[17][2] ), .C(\gbuff[18][2] ), .D(
        \gbuff[19][2] ), .S0(n1439), .S1(n1418), .Y(n56) );
  MX4X1 U523 ( .A(\gbuff[0][3] ), .B(\gbuff[1][3] ), .C(\gbuff[2][3] ), .D(
        \gbuff[3][3] ), .S0(n1440), .S1(n1419), .Y(n70) );
  MX4X1 U524 ( .A(\gbuff[16][3] ), .B(\gbuff[17][3] ), .C(\gbuff[18][3] ), .D(
        \gbuff[19][3] ), .S0(n1440), .S1(n1419), .Y(n66) );
  MX4X1 U525 ( .A(\gbuff[0][4] ), .B(\gbuff[1][4] ), .C(\gbuff[2][4] ), .D(
        \gbuff[3][4] ), .S0(n1441), .S1(n1420), .Y(n80) );
  MX4X1 U526 ( .A(\gbuff[16][4] ), .B(\gbuff[17][4] ), .C(\gbuff[18][4] ), .D(
        \gbuff[19][4] ), .S0(n1441), .S1(n1420), .Y(n76) );
  MX4X1 U527 ( .A(\gbuff[0][5] ), .B(\gbuff[1][5] ), .C(\gbuff[2][5] ), .D(
        \gbuff[3][5] ), .S0(n1441), .S1(n1420), .Y(n90) );
  MX4X1 U528 ( .A(\gbuff[16][5] ), .B(\gbuff[17][5] ), .C(\gbuff[18][5] ), .D(
        \gbuff[19][5] ), .S0(n1441), .S1(n1420), .Y(n86) );
  MX4X1 U529 ( .A(\gbuff[0][6] ), .B(\gbuff[1][6] ), .C(\gbuff[2][6] ), .D(
        \gbuff[3][6] ), .S0(n1442), .S1(n1421), .Y(n100) );
  MX4X1 U530 ( .A(\gbuff[16][6] ), .B(\gbuff[17][6] ), .C(\gbuff[18][6] ), .D(
        \gbuff[19][6] ), .S0(n1442), .S1(n1421), .Y(n96) );
  MX4X1 U531 ( .A(\gbuff[0][7] ), .B(\gbuff[1][7] ), .C(\gbuff[2][7] ), .D(
        \gbuff[3][7] ), .S0(n1443), .S1(n1421), .Y(n121) );
  MX4X1 U532 ( .A(\gbuff[16][7] ), .B(\gbuff[17][7] ), .C(\gbuff[18][7] ), .D(
        \gbuff[19][7] ), .S0(n1442), .S1(n1421), .Y(n112) );
  MX4X1 U533 ( .A(\gbuff[0][8] ), .B(\gbuff[1][8] ), .C(\gbuff[2][8] ), .D(
        \gbuff[3][8] ), .S0(n1443), .S1(n1416), .Y(n1173) );
  MX4X1 U534 ( .A(\gbuff[16][8] ), .B(\gbuff[17][8] ), .C(\gbuff[18][8] ), .D(
        \gbuff[19][8] ), .S0(n1443), .S1(n1418), .Y(n127) );
  MX4X1 U535 ( .A(\gbuff[0][9] ), .B(\gbuff[1][9] ), .C(\gbuff[2][9] ), .D(
        \gbuff[3][9] ), .S0(n1444), .S1(n1422), .Y(n1183) );
  MX4X1 U536 ( .A(\gbuff[16][9] ), .B(\gbuff[17][9] ), .C(\gbuff[18][9] ), .D(
        \gbuff[19][9] ), .S0(n1444), .S1(n1422), .Y(n1179) );
  MX4X1 U537 ( .A(\gbuff[0][10] ), .B(\gbuff[1][10] ), .C(\gbuff[2][10] ), .D(
        \gbuff[3][10] ), .S0(n1437), .S1(n1423), .Y(n1193) );
  MX4X1 U538 ( .A(\gbuff[16][10] ), .B(\gbuff[17][10] ), .C(\gbuff[18][10] ), 
        .D(\gbuff[19][10] ), .S0(n1444), .S1(n1422), .Y(n1189) );
  MX4X1 U539 ( .A(\gbuff[0][11] ), .B(\gbuff[1][11] ), .C(\gbuff[2][11] ), .D(
        \gbuff[3][11] ), .S0(n1436), .S1(n1423), .Y(n1203) );
  MX4X1 U540 ( .A(\gbuff[16][11] ), .B(\gbuff[17][11] ), .C(\gbuff[18][11] ), 
        .D(\gbuff[19][11] ), .S0(n1435), .S1(n1423), .Y(n1199) );
  MX4X1 U541 ( .A(\gbuff[0][12] ), .B(\gbuff[1][12] ), .C(\gbuff[2][12] ), .D(
        \gbuff[3][12] ), .S0(n1445), .S1(n1424), .Y(n1213) );
  MX4X1 U542 ( .A(\gbuff[16][12] ), .B(\gbuff[17][12] ), .C(\gbuff[18][12] ), 
        .D(\gbuff[19][12] ), .S0(n1437), .S1(n1423), .Y(n1209) );
  MX4X1 U543 ( .A(\gbuff[0][13] ), .B(\gbuff[1][13] ), .C(\gbuff[2][13] ), .D(
        \gbuff[3][13] ), .S0(n1445), .S1(n1424), .Y(n1223) );
  MX4X1 U544 ( .A(\gbuff[16][13] ), .B(\gbuff[17][13] ), .C(\gbuff[18][13] ), 
        .D(\gbuff[19][13] ), .S0(n1445), .S1(n1424), .Y(n1219) );
  MX4X1 U545 ( .A(\gbuff[0][14] ), .B(\gbuff[1][14] ), .C(\gbuff[2][14] ), .D(
        \gbuff[3][14] ), .S0(n1446), .S1(n1425), .Y(n1233) );
  MX4X1 U546 ( .A(\gbuff[16][14] ), .B(\gbuff[17][14] ), .C(\gbuff[18][14] ), 
        .D(\gbuff[19][14] ), .S0(n1446), .S1(n1425), .Y(n1229) );
  MX4X1 U547 ( .A(\gbuff[0][15] ), .B(\gbuff[1][15] ), .C(\gbuff[2][15] ), .D(
        \gbuff[3][15] ), .S0(n1447), .S1(n1426), .Y(n1243) );
  MX4X1 U548 ( .A(\gbuff[16][15] ), .B(\gbuff[17][15] ), .C(\gbuff[18][15] ), 
        .D(\gbuff[19][15] ), .S0(n1446), .S1(n1425), .Y(n1239) );
  MX4X1 U549 ( .A(\gbuff[0][16] ), .B(\gbuff[1][16] ), .C(\gbuff[2][16] ), .D(
        \gbuff[3][16] ), .S0(n1447), .S1(n1426), .Y(n1253) );
  MX4X1 U550 ( .A(\gbuff[16][16] ), .B(\gbuff[17][16] ), .C(\gbuff[18][16] ), 
        .D(\gbuff[19][16] ), .S0(n1447), .S1(n1426), .Y(n1249) );
  MX4X1 U551 ( .A(\gbuff[0][17] ), .B(\gbuff[1][17] ), .C(\gbuff[2][17] ), .D(
        \gbuff[3][17] ), .S0(n1434), .S1(n1427), .Y(n1263) );
  MX4X1 U552 ( .A(\gbuff[16][17] ), .B(\gbuff[17][17] ), .C(\gbuff[18][17] ), 
        .D(\gbuff[19][17] ), .S0(n1435), .S1(n1427), .Y(n1259) );
  MX4X1 U553 ( .A(\gbuff[0][18] ), .B(\gbuff[1][18] ), .C(\gbuff[2][18] ), .D(
        \gbuff[3][18] ), .S0(n1434), .S1(n1427), .Y(n1273) );
  MX4X1 U554 ( .A(\gbuff[16][18] ), .B(\gbuff[17][18] ), .C(\gbuff[18][18] ), 
        .D(\gbuff[19][18] ), .S0(n1437), .S1(n1427), .Y(n1269) );
  MX4X1 U555 ( .A(\gbuff[0][19] ), .B(\gbuff[1][19] ), .C(\gbuff[2][19] ), .D(
        \gbuff[3][19] ), .S0(n1435), .S1(n1428), .Y(n1283) );
  MX4X1 U556 ( .A(\gbuff[16][19] ), .B(\gbuff[17][19] ), .C(\gbuff[18][19] ), 
        .D(\gbuff[19][19] ), .S0(n1436), .S1(n1428), .Y(n1279) );
  MX4X1 U557 ( .A(\gbuff[0][20] ), .B(\gbuff[1][20] ), .C(\gbuff[2][20] ), .D(
        \gbuff[3][20] ), .S0(n1448), .S1(n1429), .Y(n1293) );
  MX4X1 U558 ( .A(\gbuff[16][20] ), .B(\gbuff[17][20] ), .C(\gbuff[18][20] ), 
        .D(\gbuff[19][20] ), .S0(n1437), .S1(n1428), .Y(n1289) );
  MX4X1 U559 ( .A(\gbuff[0][21] ), .B(\gbuff[1][21] ), .C(\gbuff[2][21] ), .D(
        \gbuff[3][21] ), .S0(n1448), .S1(n1429), .Y(n1303) );
  MX4X1 U560 ( .A(\gbuff[16][21] ), .B(\gbuff[17][21] ), .C(\gbuff[18][21] ), 
        .D(\gbuff[19][21] ), .S0(n1448), .S1(n1429), .Y(n1299) );
  MX4X1 U561 ( .A(\gbuff[0][22] ), .B(\gbuff[1][22] ), .C(\gbuff[2][22] ), .D(
        \gbuff[3][22] ), .S0(n1438), .S1(n1430), .Y(n1313) );
  MX4X1 U562 ( .A(\gbuff[16][22] ), .B(\gbuff[17][22] ), .C(\gbuff[18][22] ), 
        .D(\gbuff[19][22] ), .S0(N10), .S1(n1430), .Y(n1309) );
  MX4X1 U563 ( .A(\gbuff[0][23] ), .B(\gbuff[1][23] ), .C(\gbuff[2][23] ), .D(
        \gbuff[3][23] ), .S0(n1449), .S1(n1415), .Y(n1323) );
  MX4X1 U564 ( .A(\gbuff[16][23] ), .B(\gbuff[17][23] ), .C(\gbuff[18][23] ), 
        .D(\gbuff[19][23] ), .S0(N10), .S1(n1430), .Y(n1319) );
  MX4X1 U565 ( .A(\gbuff[0][24] ), .B(\gbuff[1][24] ), .C(\gbuff[2][24] ), .D(
        \gbuff[3][24] ), .S0(n1449), .S1(n1416), .Y(n1333) );
  MX4X1 U566 ( .A(\gbuff[16][24] ), .B(\gbuff[17][24] ), .C(\gbuff[18][24] ), 
        .D(\gbuff[19][24] ), .S0(n1449), .S1(n1428), .Y(n1329) );
  MX4X1 U567 ( .A(\gbuff[0][25] ), .B(\gbuff[1][25] ), .C(\gbuff[2][25] ), .D(
        \gbuff[3][25] ), .S0(n1450), .S1(n1431), .Y(n1343) );
  MX4X1 U568 ( .A(\gbuff[16][25] ), .B(\gbuff[17][25] ), .C(\gbuff[18][25] ), 
        .D(\gbuff[19][25] ), .S0(n1449), .S1(n1415), .Y(n1339) );
  MX4X1 U569 ( .A(\gbuff[0][26] ), .B(\gbuff[1][26] ), .C(\gbuff[2][26] ), .D(
        \gbuff[3][26] ), .S0(n1450), .S1(n1431), .Y(n1353) );
  MX4X1 U570 ( .A(\gbuff[16][26] ), .B(\gbuff[17][26] ), .C(\gbuff[18][26] ), 
        .D(\gbuff[19][26] ), .S0(n1450), .S1(n1431), .Y(n1349) );
  MX4X1 U571 ( .A(\gbuff[0][27] ), .B(\gbuff[1][27] ), .C(\gbuff[2][27] ), .D(
        \gbuff[3][27] ), .S0(n1451), .S1(n1432), .Y(n1363) );
  MX4X1 U572 ( .A(\gbuff[16][27] ), .B(\gbuff[17][27] ), .C(\gbuff[18][27] ), 
        .D(\gbuff[19][27] ), .S0(n1451), .S1(n1432), .Y(n1359) );
  MX4X1 U573 ( .A(\gbuff[0][28] ), .B(\gbuff[1][28] ), .C(\gbuff[2][28] ), .D(
        \gbuff[3][28] ), .S0(n1452), .S1(n1433), .Y(n1373) );
  MX4X1 U574 ( .A(\gbuff[16][28] ), .B(\gbuff[17][28] ), .C(\gbuff[18][28] ), 
        .D(\gbuff[19][28] ), .S0(n1451), .S1(n1432), .Y(n1369) );
  MX4X1 U575 ( .A(\gbuff[0][29] ), .B(\gbuff[1][29] ), .C(\gbuff[2][29] ), .D(
        \gbuff[3][29] ), .S0(n1452), .S1(n1433), .Y(n1383) );
  MX4X1 U576 ( .A(\gbuff[16][29] ), .B(\gbuff[17][29] ), .C(\gbuff[18][29] ), 
        .D(\gbuff[19][29] ), .S0(n1452), .S1(n1433), .Y(n1379) );
  MX4X1 U577 ( .A(\gbuff[0][30] ), .B(\gbuff[1][30] ), .C(\gbuff[2][30] ), .D(
        \gbuff[3][30] ), .S0(n1453), .S1(n1429), .Y(n1393) );
  MX4X1 U578 ( .A(\gbuff[16][30] ), .B(\gbuff[17][30] ), .C(\gbuff[18][30] ), 
        .D(\gbuff[19][30] ), .S0(n1453), .S1(n1425), .Y(n1389) );
  MX4X1 U579 ( .A(\gbuff[0][31] ), .B(\gbuff[1][31] ), .C(\gbuff[2][31] ), .D(
        \gbuff[3][31] ), .S0(n1453), .S1(n1424), .Y(n1403) );
  MX4X1 U580 ( .A(\gbuff[16][31] ), .B(\gbuff[17][31] ), .C(\gbuff[18][31] ), 
        .D(\gbuff[19][31] ), .S0(n1453), .S1(n1422), .Y(n1399) );
  MX4X1 U581 ( .A(\gbuff[8][0] ), .B(\gbuff[9][0] ), .C(\gbuff[10][0] ), .D(
        \gbuff[11][0] ), .S0(n1438), .S1(n1424), .Y(n38) );
  MX4X1 U582 ( .A(\gbuff[24][0] ), .B(\gbuff[25][0] ), .C(\gbuff[26][0] ), .D(
        \gbuff[27][0] ), .S0(n1438), .S1(n1425), .Y(n34) );
  MX4X1 U583 ( .A(\gbuff[8][1] ), .B(\gbuff[9][1] ), .C(\gbuff[10][1] ), .D(
        \gbuff[11][1] ), .S0(n1439), .S1(n1418), .Y(n48) );
  MX4X1 U584 ( .A(\gbuff[24][1] ), .B(\gbuff[25][1] ), .C(\gbuff[26][1] ), .D(
        \gbuff[27][1] ), .S0(n1439), .S1(n1418), .Y(n44) );
  MX4X1 U585 ( .A(\gbuff[8][2] ), .B(\gbuff[9][2] ), .C(\gbuff[10][2] ), .D(
        \gbuff[11][2] ), .S0(n1439), .S1(n1418), .Y(n58) );
  MX4X1 U586 ( .A(\gbuff[24][2] ), .B(\gbuff[25][2] ), .C(\gbuff[26][2] ), .D(
        \gbuff[27][2] ), .S0(n1439), .S1(n1418), .Y(n54) );
  MX4X1 U587 ( .A(\gbuff[8][3] ), .B(\gbuff[9][3] ), .C(\gbuff[10][3] ), .D(
        \gbuff[11][3] ), .S0(n1440), .S1(n1419), .Y(n68) );
  MX4X1 U588 ( .A(\gbuff[24][3] ), .B(\gbuff[25][3] ), .C(\gbuff[26][3] ), .D(
        \gbuff[27][3] ), .S0(n1440), .S1(n1419), .Y(n64) );
  MX4X1 U589 ( .A(\gbuff[8][4] ), .B(\gbuff[9][4] ), .C(\gbuff[10][4] ), .D(
        \gbuff[11][4] ), .S0(n1441), .S1(n1420), .Y(n78) );
  MX4X1 U590 ( .A(\gbuff[24][4] ), .B(\gbuff[25][4] ), .C(\gbuff[26][4] ), .D(
        \gbuff[27][4] ), .S0(n1440), .S1(n1419), .Y(n74) );
  MX4X1 U591 ( .A(\gbuff[8][5] ), .B(\gbuff[9][5] ), .C(\gbuff[10][5] ), .D(
        \gbuff[11][5] ), .S0(n1441), .S1(n1420), .Y(n88) );
  MX4X1 U592 ( .A(\gbuff[24][5] ), .B(\gbuff[25][5] ), .C(\gbuff[26][5] ), .D(
        \gbuff[27][5] ), .S0(n1441), .S1(n1420), .Y(n84) );
  MX4X1 U593 ( .A(\gbuff[8][6] ), .B(\gbuff[9][6] ), .C(\gbuff[10][6] ), .D(
        \gbuff[11][6] ), .S0(n1442), .S1(n1421), .Y(n98) );
  MX4X1 U594 ( .A(\gbuff[24][6] ), .B(\gbuff[25][6] ), .C(\gbuff[26][6] ), .D(
        \gbuff[27][6] ), .S0(n1442), .S1(n1421), .Y(n94) );
  MX4X1 U595 ( .A(\gbuff[8][7] ), .B(\gbuff[9][7] ), .C(\gbuff[10][7] ), .D(
        \gbuff[11][7] ), .S0(n1443), .S1(n1426), .Y(n116) );
  MX4X1 U596 ( .A(\gbuff[24][7] ), .B(\gbuff[25][7] ), .C(\gbuff[26][7] ), .D(
        \gbuff[27][7] ), .S0(n1442), .S1(n1421), .Y(n108) );
  MX4X1 U597 ( .A(\gbuff[8][8] ), .B(\gbuff[9][8] ), .C(\gbuff[10][8] ), .D(
        \gbuff[11][8] ), .S0(n1443), .S1(n1429), .Y(n1171) );
  MX4X1 U598 ( .A(\gbuff[24][8] ), .B(\gbuff[25][8] ), .C(\gbuff[26][8] ), .D(
        \gbuff[27][8] ), .S0(n1443), .S1(n1432), .Y(n125) );
  MX4X1 U599 ( .A(\gbuff[8][9] ), .B(\gbuff[9][9] ), .C(\gbuff[10][9] ), .D(
        \gbuff[11][9] ), .S0(n1444), .S1(n1422), .Y(n1181) );
  MX4X1 U600 ( .A(\gbuff[24][9] ), .B(\gbuff[25][9] ), .C(\gbuff[26][9] ), .D(
        \gbuff[27][9] ), .S0(n1443), .S1(n1433), .Y(n1177) );
  MX4X1 U601 ( .A(\gbuff[8][10] ), .B(\gbuff[9][10] ), .C(\gbuff[10][10] ), 
        .D(\gbuff[11][10] ), .S0(n1444), .S1(n1422), .Y(n1191) );
  MX4X1 U602 ( .A(\gbuff[24][10] ), .B(\gbuff[25][10] ), .C(\gbuff[26][10] ), 
        .D(\gbuff[27][10] ), .S0(n1444), .S1(n1422), .Y(n1187) );
  MX4X1 U603 ( .A(\gbuff[8][11] ), .B(\gbuff[9][11] ), .C(\gbuff[10][11] ), 
        .D(\gbuff[11][11] ), .S0(n1436), .S1(n1423), .Y(n1201) );
  MX4X1 U604 ( .A(\gbuff[24][11] ), .B(\gbuff[25][11] ), .C(\gbuff[26][11] ), 
        .D(\gbuff[27][11] ), .S0(n1436), .S1(n1423), .Y(n1197) );
  MX4X1 U605 ( .A(\gbuff[8][12] ), .B(\gbuff[9][12] ), .C(\gbuff[10][12] ), 
        .D(\gbuff[11][12] ), .S0(n1445), .S1(n1424), .Y(n1211) );
  MX4X1 U606 ( .A(\gbuff[24][12] ), .B(\gbuff[25][12] ), .C(\gbuff[26][12] ), 
        .D(\gbuff[27][12] ), .S0(n1435), .S1(n1423), .Y(n1207) );
  MX4X1 U607 ( .A(\gbuff[8][13] ), .B(\gbuff[9][13] ), .C(\gbuff[10][13] ), 
        .D(\gbuff[11][13] ), .S0(n1445), .S1(n1424), .Y(n1221) );
  MX4X1 U608 ( .A(\gbuff[24][13] ), .B(\gbuff[25][13] ), .C(\gbuff[26][13] ), 
        .D(\gbuff[27][13] ), .S0(n1445), .S1(n1424), .Y(n1217) );
  MX4X1 U609 ( .A(\gbuff[8][14] ), .B(\gbuff[9][14] ), .C(\gbuff[10][14] ), 
        .D(\gbuff[11][14] ), .S0(n1446), .S1(n1425), .Y(n1231) );
  MX4X1 U610 ( .A(\gbuff[24][14] ), .B(\gbuff[25][14] ), .C(\gbuff[26][14] ), 
        .D(\gbuff[27][14] ), .S0(n1446), .S1(n1425), .Y(n1227) );
  MX4X1 U611 ( .A(\gbuff[8][15] ), .B(\gbuff[9][15] ), .C(\gbuff[10][15] ), 
        .D(\gbuff[11][15] ), .S0(n1446), .S1(n1425), .Y(n1241) );
  MX4X1 U612 ( .A(\gbuff[24][15] ), .B(\gbuff[25][15] ), .C(\gbuff[26][15] ), 
        .D(\gbuff[27][15] ), .S0(n1446), .S1(n1425), .Y(n1237) );
  MX4X1 U613 ( .A(\gbuff[8][16] ), .B(\gbuff[9][16] ), .C(\gbuff[10][16] ), 
        .D(\gbuff[11][16] ), .S0(n1447), .S1(n1426), .Y(n1251) );
  MX4X1 U614 ( .A(\gbuff[24][16] ), .B(\gbuff[25][16] ), .C(\gbuff[26][16] ), 
        .D(\gbuff[27][16] ), .S0(n1447), .S1(n1426), .Y(n1247) );
  MX4X1 U615 ( .A(\gbuff[8][17] ), .B(\gbuff[9][17] ), .C(\gbuff[10][17] ), 
        .D(\gbuff[11][17] ), .S0(n1434), .S1(n1427), .Y(n1261) );
  MX4X1 U616 ( .A(\gbuff[24][17] ), .B(\gbuff[25][17] ), .C(\gbuff[26][17] ), 
        .D(\gbuff[27][17] ), .S0(n1447), .S1(n1426), .Y(n1257) );
  MX4X1 U617 ( .A(\gbuff[8][18] ), .B(\gbuff[9][18] ), .C(\gbuff[10][18] ), 
        .D(\gbuff[11][18] ), .S0(n1434), .S1(n1427), .Y(n1271) );
  MX4X1 U618 ( .A(\gbuff[24][18] ), .B(\gbuff[25][18] ), .C(\gbuff[26][18] ), 
        .D(\gbuff[27][18] ), .S0(n1434), .S1(n1427), .Y(n1267) );
  MX4X1 U619 ( .A(\gbuff[8][19] ), .B(\gbuff[9][19] ), .C(\gbuff[10][19] ), 
        .D(\gbuff[11][19] ), .S0(n1437), .S1(n1428), .Y(n1281) );
  MX4X1 U620 ( .A(\gbuff[24][19] ), .B(\gbuff[25][19] ), .C(\gbuff[26][19] ), 
        .D(\gbuff[27][19] ), .S0(n1437), .S1(n1428), .Y(n1277) );
  MX4X1 U621 ( .A(\gbuff[8][20] ), .B(\gbuff[9][20] ), .C(\gbuff[10][20] ), 
        .D(\gbuff[11][20] ), .S0(n1448), .S1(n1429), .Y(n1291) );
  MX4X1 U622 ( .A(\gbuff[24][20] ), .B(\gbuff[25][20] ), .C(\gbuff[26][20] ), 
        .D(\gbuff[27][20] ), .S0(n1434), .S1(n1428), .Y(n1287) );
  MX4X1 U623 ( .A(\gbuff[8][21] ), .B(\gbuff[9][21] ), .C(\gbuff[10][21] ), 
        .D(\gbuff[11][21] ), .S0(n1448), .S1(n1429), .Y(n1301) );
  MX4X1 U624 ( .A(\gbuff[24][21] ), .B(\gbuff[25][21] ), .C(\gbuff[26][21] ), 
        .D(\gbuff[27][21] ), .S0(n1448), .S1(n1429), .Y(n1297) );
  MX4X1 U625 ( .A(\gbuff[8][22] ), .B(\gbuff[9][22] ), .C(\gbuff[10][22] ), 
        .D(\gbuff[11][22] ), .S0(n1438), .S1(n1430), .Y(n1311) );
  MX4X1 U626 ( .A(\gbuff[24][22] ), .B(\gbuff[25][22] ), .C(\gbuff[26][22] ), 
        .D(\gbuff[27][22] ), .S0(n1448), .S1(n1429), .Y(n1307) );
  MX4X1 U627 ( .A(\gbuff[8][23] ), .B(\gbuff[9][23] ), .C(\gbuff[10][23] ), 
        .D(\gbuff[11][23] ), .S0(n1438), .S1(n1430), .Y(n1321) );
  MX4X1 U628 ( .A(\gbuff[24][23] ), .B(\gbuff[25][23] ), .C(\gbuff[26][23] ), 
        .D(\gbuff[27][23] ), .S0(n1438), .S1(n1430), .Y(n1317) );
  MX4X1 U629 ( .A(\gbuff[8][24] ), .B(\gbuff[9][24] ), .C(\gbuff[10][24] ), 
        .D(\gbuff[11][24] ), .S0(n1449), .S1(n1423), .Y(n1331) );
  MX4X1 U630 ( .A(\gbuff[24][24] ), .B(\gbuff[25][24] ), .C(\gbuff[26][24] ), 
        .D(\gbuff[27][24] ), .S0(n1449), .S1(n1423), .Y(n1327) );
  MX4X1 U631 ( .A(\gbuff[8][25] ), .B(\gbuff[9][25] ), .C(\gbuff[10][25] ), 
        .D(\gbuff[11][25] ), .S0(n1450), .S1(n1431), .Y(n1341) );
  MX4X1 U632 ( .A(\gbuff[24][25] ), .B(\gbuff[25][25] ), .C(\gbuff[26][25] ), 
        .D(\gbuff[27][25] ), .S0(n1449), .S1(n1417), .Y(n1337) );
  MX4X1 U633 ( .A(\gbuff[8][26] ), .B(\gbuff[9][26] ), .C(\gbuff[10][26] ), 
        .D(\gbuff[11][26] ), .S0(n1450), .S1(n1431), .Y(n1351) );
  MX4X1 U634 ( .A(\gbuff[24][26] ), .B(\gbuff[25][26] ), .C(\gbuff[26][26] ), 
        .D(\gbuff[27][26] ), .S0(n1450), .S1(n1431), .Y(n1347) );
  MX4X1 U635 ( .A(\gbuff[8][27] ), .B(\gbuff[9][27] ), .C(\gbuff[10][27] ), 
        .D(\gbuff[11][27] ), .S0(n1451), .S1(n1432), .Y(n1361) );
  MX4X1 U636 ( .A(\gbuff[24][27] ), .B(\gbuff[25][27] ), .C(\gbuff[26][27] ), 
        .D(\gbuff[27][27] ), .S0(n1451), .S1(n1432), .Y(n1357) );
  MX4X1 U637 ( .A(\gbuff[8][28] ), .B(\gbuff[9][28] ), .C(\gbuff[10][28] ), 
        .D(\gbuff[11][28] ), .S0(n1451), .S1(n1432), .Y(n1371) );
  MX4X1 U638 ( .A(\gbuff[24][28] ), .B(\gbuff[25][28] ), .C(\gbuff[26][28] ), 
        .D(\gbuff[27][28] ), .S0(n1451), .S1(n1432), .Y(n1367) );
  MX4X1 U639 ( .A(\gbuff[8][29] ), .B(\gbuff[9][29] ), .C(\gbuff[10][29] ), 
        .D(\gbuff[11][29] ), .S0(n1452), .S1(n1433), .Y(n1381) );
  MX4X1 U640 ( .A(\gbuff[24][29] ), .B(\gbuff[25][29] ), .C(\gbuff[26][29] ), 
        .D(\gbuff[27][29] ), .S0(n1452), .S1(n1433), .Y(n1377) );
  MX4X1 U641 ( .A(\gbuff[8][30] ), .B(\gbuff[9][30] ), .C(\gbuff[10][30] ), 
        .D(\gbuff[11][30] ), .S0(n1453), .S1(n1427), .Y(n1391) );
  MX4X1 U642 ( .A(\gbuff[24][30] ), .B(\gbuff[25][30] ), .C(\gbuff[26][30] ), 
        .D(\gbuff[27][30] ), .S0(n1452), .S1(n1433), .Y(n1387) );
  MX4X1 U643 ( .A(\gbuff[8][31] ), .B(\gbuff[9][31] ), .C(\gbuff[10][31] ), 
        .D(\gbuff[11][31] ), .S0(n1453), .S1(n1417), .Y(n1401) );
  MX4X1 U644 ( .A(\gbuff[24][31] ), .B(\gbuff[25][31] ), .C(\gbuff[26][31] ), 
        .D(\gbuff[27][31] ), .S0(n1453), .S1(n1422), .Y(n1397) );
  MX4X1 U645 ( .A(\gbuff[12][0] ), .B(\gbuff[13][0] ), .C(\gbuff[14][0] ), .D(
        \gbuff[15][0] ), .S0(n1438), .S1(n1426), .Y(n37) );
  MX4X1 U646 ( .A(\gbuff[12][1] ), .B(\gbuff[13][1] ), .C(\gbuff[14][1] ), .D(
        \gbuff[15][1] ), .S0(n1439), .S1(n1418), .Y(n47) );
  MX4X1 U647 ( .A(\gbuff[12][2] ), .B(\gbuff[13][2] ), .C(\gbuff[14][2] ), .D(
        \gbuff[15][2] ), .S0(n1439), .S1(n1418), .Y(n57) );
  MX4X1 U648 ( .A(\gbuff[12][3] ), .B(\gbuff[13][3] ), .C(\gbuff[14][3] ), .D(
        \gbuff[15][3] ), .S0(n1440), .S1(n1419), .Y(n67) );
  MX4X1 U649 ( .A(\gbuff[12][4] ), .B(\gbuff[13][4] ), .C(\gbuff[14][4] ), .D(
        \gbuff[15][4] ), .S0(n1441), .S1(n1420), .Y(n77) );
  MX4X1 U650 ( .A(\gbuff[12][5] ), .B(\gbuff[13][5] ), .C(\gbuff[14][5] ), .D(
        \gbuff[15][5] ), .S0(n1441), .S1(n1420), .Y(n87) );
  MX4X1 U651 ( .A(\gbuff[12][6] ), .B(\gbuff[13][6] ), .C(\gbuff[14][6] ), .D(
        \gbuff[15][6] ), .S0(n1442), .S1(n1421), .Y(n97) );
  MX4X1 U652 ( .A(\gbuff[12][7] ), .B(\gbuff[13][7] ), .C(\gbuff[14][7] ), .D(
        \gbuff[15][7] ), .S0(n1442), .S1(n1421), .Y(n114) );
  MX4X1 U653 ( .A(\gbuff[12][8] ), .B(\gbuff[13][8] ), .C(\gbuff[14][8] ), .D(
        \gbuff[15][8] ), .S0(n1443), .S1(n1419), .Y(n1170) );
  MX4X1 U654 ( .A(\gbuff[12][9] ), .B(\gbuff[13][9] ), .C(\gbuff[14][9] ), .D(
        \gbuff[15][9] ), .S0(n1444), .S1(n1422), .Y(n1180) );
  MX4X1 U655 ( .A(\gbuff[12][10] ), .B(\gbuff[13][10] ), .C(\gbuff[14][10] ), 
        .D(\gbuff[15][10] ), .S0(n1444), .S1(n1422), .Y(n1190) );
  MX4X1 U656 ( .A(\gbuff[12][11] ), .B(\gbuff[13][11] ), .C(\gbuff[14][11] ), 
        .D(\gbuff[15][11] ), .S0(n1756), .S1(n1423), .Y(n1200) );
  MX4X1 U657 ( .A(\gbuff[12][12] ), .B(\gbuff[13][12] ), .C(\gbuff[14][12] ), 
        .D(\gbuff[15][12] ), .S0(n1445), .S1(n1424), .Y(n1210) );
  MX4X1 U658 ( .A(\gbuff[12][13] ), .B(\gbuff[13][13] ), .C(\gbuff[14][13] ), 
        .D(\gbuff[15][13] ), .S0(n1445), .S1(n1424), .Y(n1220) );
  MX4X1 U659 ( .A(\gbuff[12][14] ), .B(\gbuff[13][14] ), .C(\gbuff[14][14] ), 
        .D(\gbuff[15][14] ), .S0(n1446), .S1(n1425), .Y(n1230) );
  MX4X1 U660 ( .A(\gbuff[12][15] ), .B(\gbuff[13][15] ), .C(\gbuff[14][15] ), 
        .D(\gbuff[15][15] ), .S0(n1446), .S1(n1425), .Y(n1240) );
  MX4X1 U661 ( .A(\gbuff[12][16] ), .B(\gbuff[13][16] ), .C(\gbuff[14][16] ), 
        .D(\gbuff[15][16] ), .S0(n1447), .S1(n1426), .Y(n1250) );
  MX4X1 U662 ( .A(\gbuff[12][17] ), .B(\gbuff[13][17] ), .C(\gbuff[14][17] ), 
        .D(\gbuff[15][17] ), .S0(n1436), .S1(n1427), .Y(n1260) );
  MX4X1 U663 ( .A(\gbuff[12][18] ), .B(\gbuff[13][18] ), .C(\gbuff[14][18] ), 
        .D(\gbuff[15][18] ), .S0(n1435), .S1(n1427), .Y(n1270) );
  MX4X1 U664 ( .A(\gbuff[12][19] ), .B(\gbuff[13][19] ), .C(\gbuff[14][19] ), 
        .D(\gbuff[15][19] ), .S0(n1435), .S1(n1428), .Y(n1280) );
  MX4X1 U665 ( .A(\gbuff[12][20] ), .B(\gbuff[13][20] ), .C(\gbuff[14][20] ), 
        .D(\gbuff[15][20] ), .S0(n1436), .S1(n1428), .Y(n1290) );
  MX4X1 U666 ( .A(\gbuff[12][21] ), .B(\gbuff[13][21] ), .C(\gbuff[14][21] ), 
        .D(\gbuff[15][21] ), .S0(n1448), .S1(n1429), .Y(n1300) );
  MX4X1 U667 ( .A(\gbuff[12][22] ), .B(\gbuff[13][22] ), .C(\gbuff[14][22] ), 
        .D(\gbuff[15][22] ), .S0(N10), .S1(n1430), .Y(n1310) );
  MX4X1 U668 ( .A(\gbuff[12][23] ), .B(\gbuff[13][23] ), .C(\gbuff[14][23] ), 
        .D(\gbuff[15][23] ), .S0(N10), .S1(n1430), .Y(n1320) );
  MX4X1 U669 ( .A(\gbuff[12][24] ), .B(\gbuff[13][24] ), .C(\gbuff[14][24] ), 
        .D(\gbuff[15][24] ), .S0(n1449), .S1(n1415), .Y(n1330) );
  MX4X1 U670 ( .A(\gbuff[12][25] ), .B(\gbuff[13][25] ), .C(\gbuff[14][25] ), 
        .D(\gbuff[15][25] ), .S0(n1450), .S1(n1431), .Y(n1340) );
  MX4X1 U671 ( .A(\gbuff[12][26] ), .B(\gbuff[13][26] ), .C(\gbuff[14][26] ), 
        .D(\gbuff[15][26] ), .S0(n1450), .S1(n1431), .Y(n1350) );
  MX4X1 U672 ( .A(\gbuff[12][27] ), .B(\gbuff[13][27] ), .C(\gbuff[14][27] ), 
        .D(\gbuff[15][27] ), .S0(n1451), .S1(n1432), .Y(n1360) );
  MX4X1 U673 ( .A(\gbuff[12][28] ), .B(\gbuff[13][28] ), .C(\gbuff[14][28] ), 
        .D(\gbuff[15][28] ), .S0(n1451), .S1(n1432), .Y(n1370) );
  MX4X1 U674 ( .A(\gbuff[12][29] ), .B(\gbuff[13][29] ), .C(\gbuff[14][29] ), 
        .D(\gbuff[15][29] ), .S0(n1452), .S1(n1433), .Y(n1380) );
  MX4X1 U675 ( .A(\gbuff[12][30] ), .B(\gbuff[13][30] ), .C(\gbuff[14][30] ), 
        .D(\gbuff[15][30] ), .S0(n1453), .S1(n1427), .Y(n1390) );
  MX4X1 U676 ( .A(\gbuff[12][31] ), .B(\gbuff[13][31] ), .C(\gbuff[14][31] ), 
        .D(\gbuff[15][31] ), .S0(n1453), .S1(n1430), .Y(n1400) );
  MXI2X1 U677 ( .A(n41), .B(n42), .S0(n1406), .Y(N47) );
  MXI4X1 U678 ( .A(n36), .B(n34), .C(n35), .D(n33), .S0(N13), .S1(n1412), .Y(
        n42) );
  MXI4X1 U679 ( .A(n40), .B(n38), .C(n39), .D(n37), .S0(n1408), .S1(n1413), 
        .Y(n41) );
  MX4X1 U680 ( .A(\gbuff[28][0] ), .B(\gbuff[29][0] ), .C(\gbuff[30][0] ), .D(
        \gbuff[31][0] ), .S0(n1438), .S1(n1427), .Y(n33) );
  MXI2X1 U681 ( .A(n51), .B(n52), .S0(n1407), .Y(N46) );
  MXI4X1 U682 ( .A(n46), .B(n44), .C(n45), .D(n43), .S0(n1408), .S1(n1414), 
        .Y(n52) );
  MXI4X1 U683 ( .A(n50), .B(n48), .C(n49), .D(n47), .S0(n1411), .S1(n1412), 
        .Y(n51) );
  MX4X1 U684 ( .A(\gbuff[28][1] ), .B(\gbuff[29][1] ), .C(\gbuff[30][1] ), .D(
        \gbuff[31][1] ), .S0(n1438), .S1(n1429), .Y(n43) );
  MXI2X1 U685 ( .A(n61), .B(n62), .S0(N14), .Y(N45) );
  MXI4X1 U686 ( .A(n56), .B(n54), .C(n55), .D(n53), .S0(n1408), .S1(n1413), 
        .Y(n62) );
  MXI4X1 U687 ( .A(n60), .B(n58), .C(n59), .D(n57), .S0(n1408), .S1(n1413), 
        .Y(n61) );
  MX4X1 U688 ( .A(\gbuff[28][2] ), .B(\gbuff[29][2] ), .C(\gbuff[30][2] ), .D(
        \gbuff[31][2] ), .S0(n1439), .S1(n1418), .Y(n53) );
  MXI2X1 U689 ( .A(n71), .B(n72), .S0(N14), .Y(N44) );
  MXI4X1 U690 ( .A(n66), .B(n64), .C(n65), .D(n63), .S0(n1408), .S1(n1413), 
        .Y(n72) );
  MXI4X1 U691 ( .A(n70), .B(n68), .C(n69), .D(n67), .S0(n1408), .S1(n1413), 
        .Y(n71) );
  MX4X1 U692 ( .A(\gbuff[28][3] ), .B(\gbuff[29][3] ), .C(\gbuff[30][3] ), .D(
        \gbuff[31][3] ), .S0(n1440), .S1(n1419), .Y(n63) );
  MXI2X1 U693 ( .A(n81), .B(n82), .S0(N14), .Y(N43) );
  MXI4X1 U694 ( .A(n76), .B(n74), .C(n75), .D(n73), .S0(n1408), .S1(n1413), 
        .Y(n82) );
  MXI4X1 U695 ( .A(n80), .B(n78), .C(n79), .D(n77), .S0(n1408), .S1(n1413), 
        .Y(n81) );
  MX4X1 U696 ( .A(\gbuff[28][4] ), .B(\gbuff[29][4] ), .C(\gbuff[30][4] ), .D(
        \gbuff[31][4] ), .S0(n1440), .S1(n1419), .Y(n73) );
  MXI2X1 U697 ( .A(n91), .B(n92), .S0(N14), .Y(N42) );
  MXI4X1 U698 ( .A(n86), .B(n84), .C(n85), .D(n83), .S0(n1408), .S1(n1413), 
        .Y(n92) );
  MXI4X1 U699 ( .A(n90), .B(n88), .C(n89), .D(n87), .S0(n1408), .S1(n1413), 
        .Y(n91) );
  MX4X1 U700 ( .A(\gbuff[28][5] ), .B(\gbuff[29][5] ), .C(\gbuff[30][5] ), .D(
        \gbuff[31][5] ), .S0(n1441), .S1(n1420), .Y(n83) );
  MXI2X1 U701 ( .A(n101), .B(n104), .S0(N14), .Y(N41) );
  MXI4X1 U702 ( .A(n96), .B(n94), .C(n95), .D(n93), .S0(n1408), .S1(n1413), 
        .Y(n104) );
  MXI4X1 U703 ( .A(n100), .B(n98), .C(n99), .D(n97), .S0(n1408), .S1(n1413), 
        .Y(n101) );
  MX4X1 U704 ( .A(\gbuff[28][6] ), .B(\gbuff[29][6] ), .C(\gbuff[30][6] ), .D(
        \gbuff[31][6] ), .S0(n1442), .S1(n1421), .Y(n93) );
  MXI2X1 U705 ( .A(n122), .B(n123), .S0(N14), .Y(N40) );
  MXI4X1 U706 ( .A(n112), .B(n108), .C(n110), .D(n106), .S0(n1408), .S1(n1413), 
        .Y(n123) );
  MXI4X1 U707 ( .A(n121), .B(n116), .C(n119), .D(n114), .S0(n1408), .S1(n1413), 
        .Y(n122) );
  MX4X1 U708 ( .A(\gbuff[28][7] ), .B(\gbuff[29][7] ), .C(\gbuff[30][7] ), .D(
        \gbuff[31][7] ), .S0(n1442), .S1(n1421), .Y(n106) );
  MXI2X1 U709 ( .A(n1174), .B(n1175), .S0(n1406), .Y(N39) );
  MXI4X1 U710 ( .A(n127), .B(n125), .C(n126), .D(n124), .S0(n1409), .S1(n1414), 
        .Y(n1175) );
  MXI4X1 U711 ( .A(n1173), .B(n1171), .C(n1172), .D(n1170), .S0(n1410), .S1(
        n1414), .Y(n1174) );
  MX4X1 U712 ( .A(\gbuff[28][8] ), .B(\gbuff[29][8] ), .C(\gbuff[30][8] ), .D(
        \gbuff[31][8] ), .S0(n1443), .S1(n1420), .Y(n124) );
  MXI2X1 U713 ( .A(n1184), .B(n1185), .S0(n1406), .Y(N38) );
  MXI4X1 U714 ( .A(n1179), .B(n1177), .C(n1178), .D(n1176), .S0(n1408), .S1(
        n1414), .Y(n1185) );
  MXI4X1 U715 ( .A(n1183), .B(n1181), .C(n1182), .D(n1180), .S0(n1409), .S1(
        n1414), .Y(n1184) );
  MX4X1 U716 ( .A(\gbuff[28][9] ), .B(\gbuff[29][9] ), .C(\gbuff[30][9] ), .D(
        \gbuff[31][9] ), .S0(n1443), .S1(n1416), .Y(n1176) );
  MXI2X1 U717 ( .A(n1194), .B(n1195), .S0(n1406), .Y(N37) );
  MXI4X1 U718 ( .A(n1189), .B(n1187), .C(n1188), .D(n1186), .S0(N13), .S1(
        n1414), .Y(n1195) );
  MXI4X1 U719 ( .A(n1193), .B(n1191), .C(n1192), .D(n1190), .S0(n1410), .S1(
        n1414), .Y(n1194) );
  MX4X1 U720 ( .A(\gbuff[28][10] ), .B(\gbuff[29][10] ), .C(\gbuff[30][10] ), 
        .D(\gbuff[31][10] ), .S0(n1444), .S1(n1422), .Y(n1186) );
  MXI2X1 U721 ( .A(n1204), .B(n1205), .S0(n1406), .Y(N36) );
  MXI4X1 U722 ( .A(n1199), .B(n1197), .C(n1198), .D(n1196), .S0(N13), .S1(
        n1414), .Y(n1205) );
  MXI4X1 U723 ( .A(n1203), .B(n1201), .C(n1202), .D(n1200), .S0(n1409), .S1(
        n1414), .Y(n1204) );
  MX4X1 U724 ( .A(\gbuff[28][11] ), .B(\gbuff[29][11] ), .C(\gbuff[30][11] ), 
        .D(\gbuff[31][11] ), .S0(n1436), .S1(n1423), .Y(n1196) );
  MXI2X1 U725 ( .A(n1214), .B(n1215), .S0(n1406), .Y(N35) );
  MXI4X1 U726 ( .A(n1209), .B(n1207), .C(n1208), .D(n1206), .S0(n1411), .S1(
        n1414), .Y(n1215) );
  MXI4X1 U727 ( .A(n1213), .B(n1211), .C(n1212), .D(n1210), .S0(n1411), .S1(
        n1414), .Y(n1214) );
  MX4X1 U728 ( .A(\gbuff[28][12] ), .B(\gbuff[29][12] ), .C(\gbuff[30][12] ), 
        .D(\gbuff[31][12] ), .S0(n1435), .S1(n1423), .Y(n1206) );
  MXI2X1 U729 ( .A(n1224), .B(n1225), .S0(n1406), .Y(N34) );
  MXI4X1 U730 ( .A(n1219), .B(n1217), .C(n1218), .D(n1216), .S0(N13), .S1(
        n1414), .Y(n1225) );
  MXI4X1 U731 ( .A(n1223), .B(n1221), .C(n1222), .D(n1220), .S0(n1410), .S1(
        n1414), .Y(n1224) );
  MX4X1 U732 ( .A(\gbuff[28][13] ), .B(\gbuff[29][13] ), .C(\gbuff[30][13] ), 
        .D(\gbuff[31][13] ), .S0(n1445), .S1(n1424), .Y(n1216) );
  MXI2X1 U733 ( .A(n1234), .B(n1235), .S0(n1406), .Y(N33) );
  MXI4X1 U734 ( .A(n1229), .B(n1227), .C(n1228), .D(n1226), .S0(n1409), .S1(
        n1760), .Y(n1235) );
  MXI4X1 U735 ( .A(n1233), .B(n1231), .C(n1232), .D(n1230), .S0(n1409), .S1(
        n1760), .Y(n1234) );
  MX4X1 U736 ( .A(\gbuff[28][14] ), .B(\gbuff[29][14] ), .C(\gbuff[30][14] ), 
        .D(\gbuff[31][14] ), .S0(n1445), .S1(n1424), .Y(n1226) );
  MXI2X1 U737 ( .A(n1244), .B(n1245), .S0(n1406), .Y(N32) );
  MXI4X1 U738 ( .A(n1239), .B(n1237), .C(n1238), .D(n1236), .S0(n1409), .S1(
        n1760), .Y(n1245) );
  MXI4X1 U739 ( .A(n1243), .B(n1241), .C(n1242), .D(n1240), .S0(n1409), .S1(
        n1760), .Y(n1244) );
  MX4X1 U740 ( .A(\gbuff[28][15] ), .B(\gbuff[29][15] ), .C(\gbuff[30][15] ), 
        .D(\gbuff[31][15] ), .S0(n1446), .S1(n1425), .Y(n1236) );
  MXI2X1 U741 ( .A(n1254), .B(n1255), .S0(n1406), .Y(N31) );
  MXI4X1 U742 ( .A(n1249), .B(n1247), .C(n1248), .D(n1246), .S0(n1409), .S1(
        n1760), .Y(n1255) );
  MXI4X1 U743 ( .A(n1253), .B(n1251), .C(n1252), .D(n1250), .S0(n1409), .S1(
        n1414), .Y(n1254) );
  MX4X1 U744 ( .A(\gbuff[28][16] ), .B(\gbuff[29][16] ), .C(\gbuff[30][16] ), 
        .D(\gbuff[31][16] ), .S0(n1447), .S1(n1426), .Y(n1246) );
  MXI2X1 U745 ( .A(n1264), .B(n1265), .S0(n1406), .Y(N30) );
  MXI4X1 U746 ( .A(n1259), .B(n1257), .C(n1258), .D(n1256), .S0(n1409), .S1(
        n1760), .Y(n1265) );
  MXI4X1 U747 ( .A(n1263), .B(n1261), .C(n1262), .D(n1260), .S0(n1409), .S1(
        n1414), .Y(n1264) );
  MX4X1 U748 ( .A(\gbuff[28][17] ), .B(\gbuff[29][17] ), .C(\gbuff[30][17] ), 
        .D(\gbuff[31][17] ), .S0(n1447), .S1(n1426), .Y(n1256) );
  MXI2X1 U749 ( .A(n1274), .B(n1275), .S0(n1406), .Y(N29) );
  MXI4X1 U750 ( .A(n1269), .B(n1267), .C(n1268), .D(n1266), .S0(n1409), .S1(
        n1760), .Y(n1275) );
  MXI4X1 U751 ( .A(n1273), .B(n1271), .C(n1272), .D(n1270), .S0(n1409), .S1(
        n1414), .Y(n1274) );
  MX4X1 U752 ( .A(\gbuff[28][18] ), .B(\gbuff[29][18] ), .C(\gbuff[30][18] ), 
        .D(\gbuff[31][18] ), .S0(n1437), .S1(n1427), .Y(n1266) );
  MXI2X1 U753 ( .A(n1284), .B(n1285), .S0(n1406), .Y(N28) );
  MXI4X1 U754 ( .A(n1279), .B(n1277), .C(n1278), .D(n1276), .S0(n1409), .S1(
        n1760), .Y(n1285) );
  MXI4X1 U755 ( .A(n1283), .B(n1281), .C(n1282), .D(n1280), .S0(n1409), .S1(
        n1414), .Y(n1284) );
  MX4X1 U756 ( .A(\gbuff[28][19] ), .B(\gbuff[29][19] ), .C(\gbuff[30][19] ), 
        .D(\gbuff[31][19] ), .S0(n1437), .S1(n1428), .Y(n1276) );
  MXI2X1 U757 ( .A(n1294), .B(n1295), .S0(n1407), .Y(N27) );
  MXI4X1 U758 ( .A(n1289), .B(n1287), .C(n1288), .D(n1286), .S0(n1410), .S1(
        n1412), .Y(n1295) );
  MXI4X1 U759 ( .A(n1293), .B(n1291), .C(n1292), .D(n1290), .S0(n1410), .S1(
        n1412), .Y(n1294) );
  MX4X1 U760 ( .A(\gbuff[28][20] ), .B(\gbuff[29][20] ), .C(\gbuff[30][20] ), 
        .D(\gbuff[31][20] ), .S0(n1435), .S1(n1428), .Y(n1286) );
  MXI2X1 U761 ( .A(n1304), .B(n1305), .S0(n1407), .Y(N26) );
  MXI4X1 U762 ( .A(n1299), .B(n1297), .C(n1298), .D(n1296), .S0(n1410), .S1(
        n1412), .Y(n1305) );
  MXI4X1 U763 ( .A(n1303), .B(n1301), .C(n1302), .D(n1300), .S0(n1410), .S1(
        n1412), .Y(n1304) );
  MX4X1 U764 ( .A(\gbuff[28][21] ), .B(\gbuff[29][21] ), .C(\gbuff[30][21] ), 
        .D(\gbuff[31][21] ), .S0(n1448), .S1(n1429), .Y(n1296) );
  MXI2X1 U765 ( .A(n1314), .B(n1315), .S0(n1407), .Y(N25) );
  MXI4X1 U766 ( .A(n1309), .B(n1307), .C(n1308), .D(n1306), .S0(n1410), .S1(
        n1414), .Y(n1315) );
  MXI4X1 U767 ( .A(n1313), .B(n1311), .C(n1312), .D(n1310), .S0(n1410), .S1(
        n1760), .Y(n1314) );
  MX4X1 U768 ( .A(\gbuff[28][22] ), .B(\gbuff[29][22] ), .C(\gbuff[30][22] ), 
        .D(\gbuff[31][22] ), .S0(n1448), .S1(n1429), .Y(n1306) );
  MXI2X1 U769 ( .A(n1324), .B(n1325), .S0(n1407), .Y(N24) );
  MXI4X1 U770 ( .A(n1319), .B(n1317), .C(n1318), .D(n1316), .S0(n1410), .S1(
        n1414), .Y(n1325) );
  MXI4X1 U771 ( .A(n1323), .B(n1321), .C(n1322), .D(n1320), .S0(n1410), .S1(
        N12), .Y(n1324) );
  MX4X1 U772 ( .A(\gbuff[28][23] ), .B(\gbuff[29][23] ), .C(\gbuff[30][23] ), 
        .D(\gbuff[31][23] ), .S0(N10), .S1(n1430), .Y(n1316) );
  MXI2X1 U773 ( .A(n1334), .B(n1335), .S0(n1407), .Y(N23) );
  MXI4X1 U774 ( .A(n1329), .B(n1327), .C(n1328), .D(n1326), .S0(n1410), .S1(
        n1760), .Y(n1335) );
  MXI4X1 U775 ( .A(n1333), .B(n1331), .C(n1332), .D(n1330), .S0(n1410), .S1(
        n1412), .Y(n1334) );
  MX4X1 U776 ( .A(\gbuff[28][24] ), .B(\gbuff[29][24] ), .C(\gbuff[30][24] ), 
        .D(\gbuff[31][24] ), .S0(n1449), .S1(n1426), .Y(n1326) );
  MXI2X1 U777 ( .A(n1344), .B(n1345), .S0(n1407), .Y(N22) );
  MXI4X1 U778 ( .A(n1339), .B(n1337), .C(n1338), .D(n1336), .S0(n1410), .S1(
        n1414), .Y(n1345) );
  MXI4X1 U779 ( .A(n1343), .B(n1341), .C(n1342), .D(n1340), .S0(n1410), .S1(
        n1412), .Y(n1344) );
  MX4X1 U780 ( .A(\gbuff[28][25] ), .B(\gbuff[29][25] ), .C(\gbuff[30][25] ), 
        .D(\gbuff[31][25] ), .S0(n1449), .S1(n1430), .Y(n1336) );
  MXI2X1 U781 ( .A(n1354), .B(n1355), .S0(n1407), .Y(N21) );
  MXI4X1 U782 ( .A(n1349), .B(n1347), .C(n1348), .D(n1346), .S0(n1411), .S1(
        n1412), .Y(n1355) );
  MXI4X1 U783 ( .A(n1353), .B(n1351), .C(n1352), .D(n1350), .S0(n1411), .S1(
        n1412), .Y(n1354) );
  MX4X1 U784 ( .A(\gbuff[28][26] ), .B(\gbuff[29][26] ), .C(\gbuff[30][26] ), 
        .D(\gbuff[31][26] ), .S0(n1450), .S1(n1431), .Y(n1346) );
  MXI2X1 U785 ( .A(n1364), .B(n1365), .S0(n1407), .Y(N20) );
  MXI4X1 U786 ( .A(n1359), .B(n1357), .C(n1358), .D(n1356), .S0(n1411), .S1(
        n1412), .Y(n1365) );
  MXI4X1 U787 ( .A(n1363), .B(n1361), .C(n1362), .D(n1360), .S0(n1411), .S1(
        n1412), .Y(n1364) );
  MX4X1 U788 ( .A(\gbuff[28][27] ), .B(\gbuff[29][27] ), .C(\gbuff[30][27] ), 
        .D(\gbuff[31][27] ), .S0(n1450), .S1(n1431), .Y(n1356) );
  MXI2X1 U789 ( .A(n1374), .B(n1375), .S0(n1407), .Y(N19) );
  MXI4X1 U790 ( .A(n1369), .B(n1367), .C(n1368), .D(n1366), .S0(n1411), .S1(
        n1412), .Y(n1375) );
  MXI4X1 U791 ( .A(n1373), .B(n1371), .C(n1372), .D(n1370), .S0(n1411), .S1(
        n1412), .Y(n1374) );
  MX4X1 U792 ( .A(\gbuff[28][28] ), .B(\gbuff[29][28] ), .C(\gbuff[30][28] ), 
        .D(\gbuff[31][28] ), .S0(n1451), .S1(n1432), .Y(n1366) );
  MXI2X1 U793 ( .A(n1384), .B(n1385), .S0(n1407), .Y(N18) );
  MXI4X1 U794 ( .A(n1379), .B(n1377), .C(n1378), .D(n1376), .S0(n1411), .S1(
        n1412), .Y(n1385) );
  MXI4X1 U795 ( .A(n1383), .B(n1381), .C(n1382), .D(n1380), .S0(n1411), .S1(
        n1412), .Y(n1384) );
  MX4X1 U796 ( .A(\gbuff[28][29] ), .B(\gbuff[29][29] ), .C(\gbuff[30][29] ), 
        .D(\gbuff[31][29] ), .S0(n1452), .S1(n1433), .Y(n1376) );
  MXI2X1 U797 ( .A(n1394), .B(n1395), .S0(n1407), .Y(N17) );
  MXI4X1 U798 ( .A(n1389), .B(n1387), .C(n1388), .D(n1386), .S0(n1411), .S1(
        n1412), .Y(n1395) );
  MXI4X1 U799 ( .A(n1393), .B(n1391), .C(n1392), .D(n1390), .S0(n1411), .S1(
        n1412), .Y(n1394) );
  MX4X1 U800 ( .A(\gbuff[28][30] ), .B(\gbuff[29][30] ), .C(\gbuff[30][30] ), 
        .D(\gbuff[31][30] ), .S0(n1452), .S1(n1433), .Y(n1386) );
  MXI2X1 U801 ( .A(n1404), .B(n1405), .S0(n1407), .Y(N16) );
  MXI4X1 U802 ( .A(n1399), .B(n1397), .C(n1398), .D(n1396), .S0(n1411), .S1(
        n1413), .Y(n1405) );
  MXI4X1 U803 ( .A(n1403), .B(n1401), .C(n1402), .D(n1400), .S0(n1411), .S1(
        n1412), .Y(n1404) );
  MX4X1 U804 ( .A(\gbuff[28][31] ), .B(\gbuff[29][31] ), .C(\gbuff[30][31] ), 
        .D(\gbuff[31][31] ), .S0(n1453), .S1(n1429), .Y(n1396) );
  OAI2BB2XL U805 ( .B0(n1752), .B1(n1517), .A0N(\gbuff[0][0] ), .A1N(n1754), 
        .Y(n2818) );
  OAI2BB2XL U806 ( .B0(n1753), .B1(n1515), .A0N(\gbuff[0][1] ), .A1N(n1752), 
        .Y(n2817) );
  OAI2BB2XL U807 ( .B0(n1752), .B1(n1513), .A0N(\gbuff[0][2] ), .A1N(n1752), 
        .Y(n2816) );
  OAI2BB2XL U808 ( .B0(n1752), .B1(n1511), .A0N(\gbuff[0][3] ), .A1N(n1754), 
        .Y(n2815) );
  OAI2BB2XL U809 ( .B0(n1753), .B1(n1509), .A0N(\gbuff[0][4] ), .A1N(n1754), 
        .Y(n2814) );
  OAI2BB2XL U810 ( .B0(n1752), .B1(n1507), .A0N(\gbuff[0][5] ), .A1N(n1754), 
        .Y(n2813) );
  OAI2BB2XL U811 ( .B0(n1753), .B1(n1505), .A0N(\gbuff[0][6] ), .A1N(n1754), 
        .Y(n2812) );
  OAI2BB2XL U812 ( .B0(n1752), .B1(n1503), .A0N(\gbuff[0][7] ), .A1N(n1754), 
        .Y(n2811) );
  OAI2BB2XL U813 ( .B0(n1753), .B1(n1501), .A0N(\gbuff[0][8] ), .A1N(n1754), 
        .Y(n2810) );
  OAI2BB2XL U814 ( .B0(n1752), .B1(n1499), .A0N(\gbuff[0][9] ), .A1N(n1754), 
        .Y(n2809) );
  OAI2BB2XL U815 ( .B0(n1753), .B1(n1497), .A0N(\gbuff[0][10] ), .A1N(n1754), 
        .Y(n2808) );
  OAI2BB2XL U816 ( .B0(n1752), .B1(n1495), .A0N(\gbuff[0][11] ), .A1N(n1754), 
        .Y(n2807) );
  OAI2BB2XL U817 ( .B0(n1753), .B1(n1493), .A0N(\gbuff[0][12] ), .A1N(n1754), 
        .Y(n2806) );
  OAI2BB2XL U818 ( .B0(n1752), .B1(n1491), .A0N(\gbuff[0][13] ), .A1N(n1754), 
        .Y(n2805) );
  OAI2BB2XL U819 ( .B0(n1752), .B1(n1489), .A0N(\gbuff[0][14] ), .A1N(n1754), 
        .Y(n2804) );
  OAI2BB2XL U820 ( .B0(n1752), .B1(n1487), .A0N(\gbuff[0][15] ), .A1N(n1753), 
        .Y(n2803) );
  OAI2BB2XL U821 ( .B0(n1752), .B1(n1485), .A0N(\gbuff[0][16] ), .A1N(n1754), 
        .Y(n2802) );
  OAI2BB2XL U822 ( .B0(n1752), .B1(n1483), .A0N(\gbuff[0][17] ), .A1N(n1753), 
        .Y(n2801) );
  OAI2BB2XL U823 ( .B0(n1752), .B1(n1481), .A0N(\gbuff[0][18] ), .A1N(n1753), 
        .Y(n2800) );
  OAI2BB2XL U824 ( .B0(n1752), .B1(n1479), .A0N(\gbuff[0][19] ), .A1N(n1753), 
        .Y(n2799) );
  OAI2BB2XL U825 ( .B0(n1752), .B1(n1477), .A0N(\gbuff[0][20] ), .A1N(n1753), 
        .Y(n2798) );
  OAI2BB2XL U826 ( .B0(n1752), .B1(n1475), .A0N(\gbuff[0][21] ), .A1N(n1753), 
        .Y(n2797) );
  OAI2BB2XL U827 ( .B0(n1752), .B1(n1473), .A0N(\gbuff[0][22] ), .A1N(n1754), 
        .Y(n2796) );
  OAI2BB2XL U828 ( .B0(n1753), .B1(n1471), .A0N(\gbuff[0][23] ), .A1N(n1753), 
        .Y(n2795) );
  OAI2BB2XL U829 ( .B0(n1752), .B1(n1469), .A0N(\gbuff[0][24] ), .A1N(n1754), 
        .Y(n2794) );
  OAI2BB2XL U830 ( .B0(n1753), .B1(n1467), .A0N(\gbuff[0][25] ), .A1N(n1754), 
        .Y(n2793) );
  OAI2BB2XL U831 ( .B0(n1753), .B1(n1465), .A0N(\gbuff[0][26] ), .A1N(n1754), 
        .Y(n2792) );
  OAI2BB2XL U832 ( .B0(n1753), .B1(n1463), .A0N(\gbuff[0][27] ), .A1N(n1754), 
        .Y(n2791) );
  OAI2BB2XL U833 ( .B0(n1753), .B1(n1461), .A0N(\gbuff[0][28] ), .A1N(n1754), 
        .Y(n2790) );
  OAI2BB2XL U834 ( .B0(n1753), .B1(n1459), .A0N(\gbuff[0][29] ), .A1N(n1754), 
        .Y(n2789) );
  OAI2BB2XL U835 ( .B0(n1753), .B1(n1457), .A0N(\gbuff[0][30] ), .A1N(n1754), 
        .Y(n2788) );
  OAI2BB2XL U836 ( .B0(n1753), .B1(n1455), .A0N(\gbuff[0][31] ), .A1N(n1752), 
        .Y(n2787) );
  OAI2BB2XL U837 ( .B0(n1793), .B1(n1749), .A0N(\gbuff[1][0] ), .A1N(n1751), 
        .Y(n2786) );
  OAI2BB2XL U838 ( .B0(n1792), .B1(n1749), .A0N(\gbuff[1][1] ), .A1N(n1751), 
        .Y(n2785) );
  OAI2BB2XL U839 ( .B0(n1791), .B1(n1749), .A0N(\gbuff[1][2] ), .A1N(n1749), 
        .Y(n2784) );
  OAI2BB2XL U840 ( .B0(n1790), .B1(n1749), .A0N(\gbuff[1][3] ), .A1N(n1751), 
        .Y(n2783) );
  OAI2BB2XL U841 ( .B0(n1789), .B1(n1749), .A0N(\gbuff[1][4] ), .A1N(n1751), 
        .Y(n2782) );
  OAI2BB2XL U842 ( .B0(n1788), .B1(n1749), .A0N(\gbuff[1][5] ), .A1N(n1751), 
        .Y(n2781) );
  OAI2BB2XL U843 ( .B0(n1787), .B1(n1749), .A0N(\gbuff[1][6] ), .A1N(n1751), 
        .Y(n2780) );
  OAI2BB2XL U844 ( .B0(n1786), .B1(n1749), .A0N(\gbuff[1][7] ), .A1N(n1751), 
        .Y(n2779) );
  OAI2BB2XL U845 ( .B0(n1785), .B1(n1749), .A0N(\gbuff[1][8] ), .A1N(n1751), 
        .Y(n2778) );
  OAI2BB2XL U846 ( .B0(n1784), .B1(n1749), .A0N(\gbuff[1][9] ), .A1N(n1751), 
        .Y(n2777) );
  OAI2BB2XL U847 ( .B0(n1783), .B1(n1749), .A0N(\gbuff[1][10] ), .A1N(n1751), 
        .Y(n2776) );
  OAI2BB2XL U848 ( .B0(n1782), .B1(n1749), .A0N(\gbuff[1][11] ), .A1N(n1751), 
        .Y(n2775) );
  OAI2BB2XL U849 ( .B0(n1781), .B1(n1749), .A0N(\gbuff[1][12] ), .A1N(n1751), 
        .Y(n2774) );
  OAI2BB2XL U850 ( .B0(n1780), .B1(n1749), .A0N(\gbuff[1][13] ), .A1N(n1751), 
        .Y(n2773) );
  OAI2BB2XL U851 ( .B0(n1779), .B1(n1750), .A0N(\gbuff[1][14] ), .A1N(n1751), 
        .Y(n2772) );
  OAI2BB2XL U852 ( .B0(n1778), .B1(n1749), .A0N(\gbuff[1][15] ), .A1N(n1750), 
        .Y(n2771) );
  OAI2BB2XL U853 ( .B0(n1777), .B1(n1750), .A0N(\gbuff[1][16] ), .A1N(n1751), 
        .Y(n2770) );
  OAI2BB2XL U854 ( .B0(n1776), .B1(n1749), .A0N(\gbuff[1][17] ), .A1N(n1750), 
        .Y(n2769) );
  OAI2BB2XL U855 ( .B0(n1775), .B1(n1750), .A0N(\gbuff[1][18] ), .A1N(n1750), 
        .Y(n2768) );
  OAI2BB2XL U856 ( .B0(n1774), .B1(n1749), .A0N(\gbuff[1][19] ), .A1N(n1750), 
        .Y(n2767) );
  OAI2BB2XL U857 ( .B0(n1773), .B1(n1750), .A0N(\gbuff[1][20] ), .A1N(n1750), 
        .Y(n2766) );
  OAI2BB2XL U858 ( .B0(n1772), .B1(n1749), .A0N(\gbuff[1][21] ), .A1N(n1750), 
        .Y(n2765) );
  OAI2BB2XL U859 ( .B0(n1771), .B1(n1750), .A0N(\gbuff[1][22] ), .A1N(n1751), 
        .Y(n2764) );
  OAI2BB2XL U860 ( .B0(n1770), .B1(n1750), .A0N(\gbuff[1][23] ), .A1N(n1750), 
        .Y(n2763) );
  OAI2BB2XL U861 ( .B0(n1769), .B1(n1749), .A0N(\gbuff[1][24] ), .A1N(n1751), 
        .Y(n2762) );
  OAI2BB2XL U862 ( .B0(n1768), .B1(n1750), .A0N(\gbuff[1][25] ), .A1N(n1751), 
        .Y(n2761) );
  OAI2BB2XL U863 ( .B0(n1767), .B1(n1750), .A0N(\gbuff[1][26] ), .A1N(n1751), 
        .Y(n2760) );
  OAI2BB2XL U864 ( .B0(n1766), .B1(n1750), .A0N(\gbuff[1][27] ), .A1N(n1751), 
        .Y(n2759) );
  OAI2BB2XL U865 ( .B0(n1765), .B1(n1750), .A0N(\gbuff[1][28] ), .A1N(n1751), 
        .Y(n2758) );
  OAI2BB2XL U866 ( .B0(n1764), .B1(n1750), .A0N(\gbuff[1][29] ), .A1N(n1751), 
        .Y(n2757) );
  OAI2BB2XL U867 ( .B0(n1763), .B1(n1750), .A0N(\gbuff[1][30] ), .A1N(n1750), 
        .Y(n2756) );
  OAI2BB2XL U868 ( .B0(n1762), .B1(n1750), .A0N(\gbuff[1][31] ), .A1N(n1749), 
        .Y(n2755) );
  OAI2BB2XL U869 ( .B0(n1793), .B1(n1746), .A0N(\gbuff[2][0] ), .A1N(n1748), 
        .Y(n2754) );
  OAI2BB2XL U870 ( .B0(n1792), .B1(n1746), .A0N(\gbuff[2][1] ), .A1N(n1748), 
        .Y(n2753) );
  OAI2BB2XL U871 ( .B0(n1791), .B1(n1746), .A0N(\gbuff[2][2] ), .A1N(n1746), 
        .Y(n2752) );
  OAI2BB2XL U872 ( .B0(n1790), .B1(n1746), .A0N(\gbuff[2][3] ), .A1N(n1748), 
        .Y(n2751) );
  OAI2BB2XL U873 ( .B0(n1789), .B1(n1746), .A0N(\gbuff[2][4] ), .A1N(n1748), 
        .Y(n2750) );
  OAI2BB2XL U874 ( .B0(n1788), .B1(n1746), .A0N(\gbuff[2][5] ), .A1N(n1748), 
        .Y(n2749) );
  OAI2BB2XL U875 ( .B0(n1787), .B1(n1746), .A0N(\gbuff[2][6] ), .A1N(n1748), 
        .Y(n2748) );
  OAI2BB2XL U876 ( .B0(n1786), .B1(n1746), .A0N(\gbuff[2][7] ), .A1N(n1748), 
        .Y(n2747) );
  OAI2BB2XL U877 ( .B0(n1785), .B1(n1746), .A0N(\gbuff[2][8] ), .A1N(n1748), 
        .Y(n2746) );
  OAI2BB2XL U878 ( .B0(n1784), .B1(n1746), .A0N(\gbuff[2][9] ), .A1N(n1748), 
        .Y(n2745) );
  OAI2BB2XL U879 ( .B0(n1783), .B1(n1746), .A0N(\gbuff[2][10] ), .A1N(n1748), 
        .Y(n2744) );
  OAI2BB2XL U880 ( .B0(n1782), .B1(n1746), .A0N(\gbuff[2][11] ), .A1N(n1748), 
        .Y(n2743) );
  OAI2BB2XL U881 ( .B0(n1781), .B1(n1746), .A0N(\gbuff[2][12] ), .A1N(n1748), 
        .Y(n2742) );
  OAI2BB2XL U882 ( .B0(n1780), .B1(n1746), .A0N(\gbuff[2][13] ), .A1N(n1748), 
        .Y(n2741) );
  OAI2BB2XL U883 ( .B0(n1779), .B1(n1747), .A0N(\gbuff[2][14] ), .A1N(n1748), 
        .Y(n2740) );
  OAI2BB2XL U884 ( .B0(n1778), .B1(n1746), .A0N(\gbuff[2][15] ), .A1N(n1747), 
        .Y(n2739) );
  OAI2BB2XL U885 ( .B0(n1777), .B1(n1747), .A0N(\gbuff[2][16] ), .A1N(n1748), 
        .Y(n2738) );
  OAI2BB2XL U886 ( .B0(n1776), .B1(n1746), .A0N(\gbuff[2][17] ), .A1N(n1747), 
        .Y(n2737) );
  OAI2BB2XL U887 ( .B0(n1775), .B1(n1747), .A0N(\gbuff[2][18] ), .A1N(n1747), 
        .Y(n2736) );
  OAI2BB2XL U888 ( .B0(n1774), .B1(n1746), .A0N(\gbuff[2][19] ), .A1N(n1747), 
        .Y(n2735) );
  OAI2BB2XL U889 ( .B0(n1773), .B1(n1747), .A0N(\gbuff[2][20] ), .A1N(n1747), 
        .Y(n2734) );
  OAI2BB2XL U890 ( .B0(n1772), .B1(n1746), .A0N(\gbuff[2][21] ), .A1N(n1747), 
        .Y(n2733) );
  OAI2BB2XL U891 ( .B0(n1771), .B1(n1747), .A0N(\gbuff[2][22] ), .A1N(n1748), 
        .Y(n2732) );
  OAI2BB2XL U892 ( .B0(n1770), .B1(n1747), .A0N(\gbuff[2][23] ), .A1N(n1747), 
        .Y(n2731) );
  OAI2BB2XL U893 ( .B0(n1769), .B1(n1746), .A0N(\gbuff[2][24] ), .A1N(n1748), 
        .Y(n2730) );
  OAI2BB2XL U894 ( .B0(n1768), .B1(n1747), .A0N(\gbuff[2][25] ), .A1N(n1748), 
        .Y(n2729) );
  OAI2BB2XL U895 ( .B0(n1767), .B1(n1747), .A0N(\gbuff[2][26] ), .A1N(n1748), 
        .Y(n2728) );
  OAI2BB2XL U896 ( .B0(n1766), .B1(n1747), .A0N(\gbuff[2][27] ), .A1N(n1748), 
        .Y(n2727) );
  OAI2BB2XL U897 ( .B0(n1765), .B1(n1747), .A0N(\gbuff[2][28] ), .A1N(n1748), 
        .Y(n2726) );
  OAI2BB2XL U898 ( .B0(n1764), .B1(n1747), .A0N(\gbuff[2][29] ), .A1N(n1748), 
        .Y(n2725) );
  OAI2BB2XL U899 ( .B0(n1763), .B1(n1747), .A0N(\gbuff[2][30] ), .A1N(n1747), 
        .Y(n2724) );
  OAI2BB2XL U900 ( .B0(n1762), .B1(n1747), .A0N(\gbuff[2][31] ), .A1N(n1746), 
        .Y(n2723) );
  OAI2BB2XL U901 ( .B0(n1793), .B1(n1743), .A0N(\gbuff[3][0] ), .A1N(n1745), 
        .Y(n2722) );
  OAI2BB2XL U902 ( .B0(n1792), .B1(n1743), .A0N(\gbuff[3][1] ), .A1N(n1745), 
        .Y(n2721) );
  OAI2BB2XL U903 ( .B0(n1791), .B1(n1743), .A0N(\gbuff[3][2] ), .A1N(n1743), 
        .Y(n2720) );
  OAI2BB2XL U904 ( .B0(n1790), .B1(n1743), .A0N(\gbuff[3][3] ), .A1N(n1745), 
        .Y(n2719) );
  OAI2BB2XL U905 ( .B0(n1789), .B1(n1743), .A0N(\gbuff[3][4] ), .A1N(n1745), 
        .Y(n2718) );
  OAI2BB2XL U906 ( .B0(n1788), .B1(n1743), .A0N(\gbuff[3][5] ), .A1N(n1745), 
        .Y(n2717) );
  OAI2BB2XL U907 ( .B0(n1787), .B1(n1743), .A0N(\gbuff[3][6] ), .A1N(n1745), 
        .Y(n2716) );
  OAI2BB2XL U908 ( .B0(n1786), .B1(n1743), .A0N(\gbuff[3][7] ), .A1N(n1745), 
        .Y(n2715) );
  OAI2BB2XL U909 ( .B0(n1785), .B1(n1743), .A0N(\gbuff[3][8] ), .A1N(n1745), 
        .Y(n2714) );
  OAI2BB2XL U910 ( .B0(n1784), .B1(n1743), .A0N(\gbuff[3][9] ), .A1N(n1745), 
        .Y(n2713) );
  OAI2BB2XL U911 ( .B0(n1783), .B1(n1743), .A0N(\gbuff[3][10] ), .A1N(n1745), 
        .Y(n2712) );
  OAI2BB2XL U912 ( .B0(n1782), .B1(n1743), .A0N(\gbuff[3][11] ), .A1N(n1745), 
        .Y(n2711) );
  OAI2BB2XL U913 ( .B0(n1781), .B1(n1743), .A0N(\gbuff[3][12] ), .A1N(n1745), 
        .Y(n2710) );
  OAI2BB2XL U914 ( .B0(n1780), .B1(n1743), .A0N(\gbuff[3][13] ), .A1N(n1745), 
        .Y(n2709) );
  OAI2BB2XL U915 ( .B0(n1779), .B1(n1744), .A0N(\gbuff[3][14] ), .A1N(n1745), 
        .Y(n2708) );
  OAI2BB2XL U916 ( .B0(n1778), .B1(n1743), .A0N(\gbuff[3][15] ), .A1N(n1744), 
        .Y(n2707) );
  OAI2BB2XL U917 ( .B0(n1777), .B1(n1744), .A0N(\gbuff[3][16] ), .A1N(n1745), 
        .Y(n2706) );
  OAI2BB2XL U918 ( .B0(n1776), .B1(n1743), .A0N(\gbuff[3][17] ), .A1N(n1744), 
        .Y(n2705) );
  OAI2BB2XL U919 ( .B0(n1775), .B1(n1744), .A0N(\gbuff[3][18] ), .A1N(n1744), 
        .Y(n2704) );
  OAI2BB2XL U920 ( .B0(n1774), .B1(n1743), .A0N(\gbuff[3][19] ), .A1N(n1744), 
        .Y(n2703) );
  OAI2BB2XL U921 ( .B0(n1773), .B1(n1744), .A0N(\gbuff[3][20] ), .A1N(n1744), 
        .Y(n2702) );
  OAI2BB2XL U922 ( .B0(n1772), .B1(n1743), .A0N(\gbuff[3][21] ), .A1N(n1744), 
        .Y(n2701) );
  OAI2BB2XL U923 ( .B0(n1771), .B1(n1744), .A0N(\gbuff[3][22] ), .A1N(n1745), 
        .Y(n2700) );
  OAI2BB2XL U924 ( .B0(n1770), .B1(n1744), .A0N(\gbuff[3][23] ), .A1N(n1744), 
        .Y(n2699) );
  OAI2BB2XL U925 ( .B0(n1769), .B1(n1743), .A0N(\gbuff[3][24] ), .A1N(n1745), 
        .Y(n2698) );
  OAI2BB2XL U926 ( .B0(n1768), .B1(n1744), .A0N(\gbuff[3][25] ), .A1N(n1745), 
        .Y(n2697) );
  OAI2BB2XL U927 ( .B0(n1767), .B1(n1744), .A0N(\gbuff[3][26] ), .A1N(n1745), 
        .Y(n2696) );
  OAI2BB2XL U928 ( .B0(n1766), .B1(n1744), .A0N(\gbuff[3][27] ), .A1N(n1745), 
        .Y(n2695) );
  OAI2BB2XL U929 ( .B0(n1765), .B1(n1744), .A0N(\gbuff[3][28] ), .A1N(n1745), 
        .Y(n2694) );
  OAI2BB2XL U930 ( .B0(n1764), .B1(n1744), .A0N(\gbuff[3][29] ), .A1N(n1745), 
        .Y(n2693) );
  OAI2BB2XL U931 ( .B0(n1763), .B1(n1744), .A0N(\gbuff[3][30] ), .A1N(n1744), 
        .Y(n2692) );
  OAI2BB2XL U932 ( .B0(n1762), .B1(n1744), .A0N(\gbuff[3][31] ), .A1N(n1743), 
        .Y(n2691) );
  OAI2BB2XL U933 ( .B0(n1793), .B1(n1741), .A0N(\gbuff[4][0] ), .A1N(n1741), 
        .Y(n2690) );
  OAI2BB2XL U934 ( .B0(n1792), .B1(n1740), .A0N(\gbuff[4][1] ), .A1N(n1740), 
        .Y(n2689) );
  OAI2BB2XL U935 ( .B0(n1791), .B1(n1740), .A0N(\gbuff[4][2] ), .A1N(n1741), 
        .Y(n2688) );
  OAI2BB2XL U936 ( .B0(n1790), .B1(n1740), .A0N(\gbuff[4][3] ), .A1N(n1742), 
        .Y(n2687) );
  OAI2BB2XL U937 ( .B0(n1789), .B1(n1740), .A0N(\gbuff[4][4] ), .A1N(n1740), 
        .Y(n2686) );
  OAI2BB2XL U938 ( .B0(n1788), .B1(n1740), .A0N(\gbuff[4][5] ), .A1N(n1742), 
        .Y(n2685) );
  OAI2BB2XL U939 ( .B0(n1787), .B1(n1740), .A0N(\gbuff[4][6] ), .A1N(n1742), 
        .Y(n2684) );
  OAI2BB2XL U940 ( .B0(n1786), .B1(n1740), .A0N(\gbuff[4][7] ), .A1N(n1742), 
        .Y(n2683) );
  OAI2BB2XL U941 ( .B0(n1785), .B1(n1740), .A0N(\gbuff[4][8] ), .A1N(n1742), 
        .Y(n2682) );
  OAI2BB2XL U942 ( .B0(n1784), .B1(n1740), .A0N(\gbuff[4][9] ), .A1N(n1742), 
        .Y(n2681) );
  OAI2BB2XL U943 ( .B0(n1783), .B1(n1740), .A0N(\gbuff[4][10] ), .A1N(n1742), 
        .Y(n2680) );
  OAI2BB2XL U944 ( .B0(n1782), .B1(n1740), .A0N(\gbuff[4][11] ), .A1N(n1742), 
        .Y(n2679) );
  OAI2BB2XL U945 ( .B0(n1781), .B1(n1740), .A0N(\gbuff[4][12] ), .A1N(n1742), 
        .Y(n2678) );
  OAI2BB2XL U946 ( .B0(n1780), .B1(n1741), .A0N(\gbuff[4][13] ), .A1N(n1742), 
        .Y(n2677) );
  OAI2BB2XL U947 ( .B0(n1779), .B1(n1741), .A0N(\gbuff[4][14] ), .A1N(n1742), 
        .Y(n2676) );
  OAI2BB2XL U948 ( .B0(n1778), .B1(n1741), .A0N(\gbuff[4][15] ), .A1N(n1741), 
        .Y(n2675) );
  OAI2BB2XL U949 ( .B0(n1777), .B1(n1741), .A0N(\gbuff[4][16] ), .A1N(n1742), 
        .Y(n2674) );
  OAI2BB2XL U950 ( .B0(n1776), .B1(n1741), .A0N(\gbuff[4][17] ), .A1N(n1740), 
        .Y(n2673) );
  OAI2BB2XL U951 ( .B0(n1775), .B1(n1741), .A0N(\gbuff[4][18] ), .A1N(n1742), 
        .Y(n2672) );
  OAI2BB2XL U952 ( .B0(n1774), .B1(n1741), .A0N(\gbuff[4][19] ), .A1N(n1741), 
        .Y(n2671) );
  OAI2BB2XL U953 ( .B0(n1773), .B1(n1741), .A0N(\gbuff[4][20] ), .A1N(n1740), 
        .Y(n2670) );
  OAI2BB2XL U954 ( .B0(n1772), .B1(n1741), .A0N(\gbuff[4][21] ), .A1N(n1742), 
        .Y(n2669) );
  OAI2BB2XL U955 ( .B0(n1771), .B1(n1741), .A0N(\gbuff[4][22] ), .A1N(n1742), 
        .Y(n2668) );
  OAI2BB2XL U956 ( .B0(n1770), .B1(n1741), .A0N(\gbuff[4][23] ), .A1N(n1742), 
        .Y(n2667) );
  OAI2BB2XL U957 ( .B0(n1769), .B1(n1741), .A0N(\gbuff[4][24] ), .A1N(n1742), 
        .Y(n2666) );
  OAI2BB2XL U958 ( .B0(n1768), .B1(n1740), .A0N(\gbuff[4][25] ), .A1N(n1742), 
        .Y(n2665) );
  OAI2BB2XL U959 ( .B0(n1767), .B1(n1741), .A0N(\gbuff[4][26] ), .A1N(n1742), 
        .Y(n2664) );
  OAI2BB2XL U960 ( .B0(n1766), .B1(n1740), .A0N(\gbuff[4][27] ), .A1N(n1742), 
        .Y(n2663) );
  OAI2BB2XL U961 ( .B0(n1765), .B1(n1741), .A0N(\gbuff[4][28] ), .A1N(n1742), 
        .Y(n2662) );
  OAI2BB2XL U962 ( .B0(n1764), .B1(n1740), .A0N(\gbuff[4][29] ), .A1N(n1742), 
        .Y(n2661) );
  OAI2BB2XL U963 ( .B0(n1763), .B1(n1741), .A0N(\gbuff[4][30] ), .A1N(n1741), 
        .Y(n2660) );
  OAI2BB2XL U964 ( .B0(n1762), .B1(n1740), .A0N(\gbuff[4][31] ), .A1N(n1740), 
        .Y(n2659) );
  OAI2BB2XL U965 ( .B0(n1793), .B1(n1737), .A0N(\gbuff[5][0] ), .A1N(n1739), 
        .Y(n2658) );
  OAI2BB2XL U966 ( .B0(n1792), .B1(n1737), .A0N(\gbuff[5][1] ), .A1N(n1739), 
        .Y(n2657) );
  OAI2BB2XL U967 ( .B0(n1791), .B1(n1737), .A0N(\gbuff[5][2] ), .A1N(n1737), 
        .Y(n2656) );
  OAI2BB2XL U968 ( .B0(n1790), .B1(n1737), .A0N(\gbuff[5][3] ), .A1N(n1739), 
        .Y(n2655) );
  OAI2BB2XL U969 ( .B0(n1789), .B1(n1737), .A0N(\gbuff[5][4] ), .A1N(n1739), 
        .Y(n2654) );
  OAI2BB2XL U970 ( .B0(n1788), .B1(n1737), .A0N(\gbuff[5][5] ), .A1N(n1739), 
        .Y(n2653) );
  OAI2BB2XL U971 ( .B0(n1787), .B1(n1737), .A0N(\gbuff[5][6] ), .A1N(n1739), 
        .Y(n2652) );
  OAI2BB2XL U972 ( .B0(n1786), .B1(n1737), .A0N(\gbuff[5][7] ), .A1N(n1739), 
        .Y(n2651) );
  OAI2BB2XL U973 ( .B0(n1785), .B1(n1737), .A0N(\gbuff[5][8] ), .A1N(n1739), 
        .Y(n2650) );
  OAI2BB2XL U974 ( .B0(n1784), .B1(n1737), .A0N(\gbuff[5][9] ), .A1N(n1739), 
        .Y(n2649) );
  OAI2BB2XL U975 ( .B0(n1783), .B1(n1737), .A0N(\gbuff[5][10] ), .A1N(n1739), 
        .Y(n2648) );
  OAI2BB2XL U976 ( .B0(n1782), .B1(n1737), .A0N(\gbuff[5][11] ), .A1N(n1739), 
        .Y(n2647) );
  OAI2BB2XL U977 ( .B0(n1781), .B1(n1737), .A0N(\gbuff[5][12] ), .A1N(n1739), 
        .Y(n2646) );
  OAI2BB2XL U978 ( .B0(n1780), .B1(n1737), .A0N(\gbuff[5][13] ), .A1N(n1739), 
        .Y(n2645) );
  OAI2BB2XL U979 ( .B0(n1779), .B1(n1738), .A0N(\gbuff[5][14] ), .A1N(n1739), 
        .Y(n2644) );
  OAI2BB2XL U980 ( .B0(n1778), .B1(n1737), .A0N(\gbuff[5][15] ), .A1N(n1738), 
        .Y(n2643) );
  OAI2BB2XL U981 ( .B0(n1777), .B1(n1738), .A0N(\gbuff[5][16] ), .A1N(n1739), 
        .Y(n2642) );
  OAI2BB2XL U982 ( .B0(n1776), .B1(n1737), .A0N(\gbuff[5][17] ), .A1N(n1738), 
        .Y(n2641) );
  OAI2BB2XL U983 ( .B0(n1775), .B1(n1738), .A0N(\gbuff[5][18] ), .A1N(n1738), 
        .Y(n2640) );
  OAI2BB2XL U984 ( .B0(n1774), .B1(n1737), .A0N(\gbuff[5][19] ), .A1N(n1738), 
        .Y(n2639) );
  OAI2BB2XL U985 ( .B0(n1773), .B1(n1738), .A0N(\gbuff[5][20] ), .A1N(n1738), 
        .Y(n2638) );
  OAI2BB2XL U986 ( .B0(n1772), .B1(n1737), .A0N(\gbuff[5][21] ), .A1N(n1738), 
        .Y(n2637) );
  OAI2BB2XL U987 ( .B0(n1771), .B1(n1738), .A0N(\gbuff[5][22] ), .A1N(n1739), 
        .Y(n2636) );
  OAI2BB2XL U988 ( .B0(n1770), .B1(n1738), .A0N(\gbuff[5][23] ), .A1N(n1738), 
        .Y(n2635) );
  OAI2BB2XL U989 ( .B0(n1769), .B1(n6), .A0N(\gbuff[5][24] ), .A1N(n1739), .Y(
        n2634) );
  OAI2BB2XL U990 ( .B0(n1768), .B1(n1738), .A0N(\gbuff[5][25] ), .A1N(n1739), 
        .Y(n2633) );
  OAI2BB2XL U991 ( .B0(n1767), .B1(n1738), .A0N(\gbuff[5][26] ), .A1N(n1739), 
        .Y(n2632) );
  OAI2BB2XL U992 ( .B0(n1766), .B1(n1738), .A0N(\gbuff[5][27] ), .A1N(n1739), 
        .Y(n2631) );
  OAI2BB2XL U993 ( .B0(n1765), .B1(n1738), .A0N(\gbuff[5][28] ), .A1N(n1739), 
        .Y(n2630) );
  OAI2BB2XL U994 ( .B0(n1764), .B1(n1738), .A0N(\gbuff[5][29] ), .A1N(n1739), 
        .Y(n2629) );
  OAI2BB2XL U995 ( .B0(n1763), .B1(n1738), .A0N(\gbuff[5][30] ), .A1N(n6), .Y(
        n2628) );
  OAI2BB2XL U996 ( .B0(n1762), .B1(n1738), .A0N(\gbuff[5][31] ), .A1N(n1737), 
        .Y(n2627) );
  OAI2BB2XL U997 ( .B0(n1517), .B1(n1734), .A0N(\gbuff[6][0] ), .A1N(n1736), 
        .Y(n2626) );
  OAI2BB2XL U998 ( .B0(n1515), .B1(n1734), .A0N(\gbuff[6][1] ), .A1N(n7), .Y(
        n2625) );
  OAI2BB2XL U999 ( .B0(n1513), .B1(n1734), .A0N(\gbuff[6][2] ), .A1N(n1734), 
        .Y(n2624) );
  OAI2BB2XL U1000 ( .B0(n1511), .B1(n1734), .A0N(\gbuff[6][3] ), .A1N(n1736), 
        .Y(n2623) );
  OAI2BB2XL U1001 ( .B0(n1509), .B1(n1734), .A0N(\gbuff[6][4] ), .A1N(n1736), 
        .Y(n2622) );
  OAI2BB2XL U1002 ( .B0(n1507), .B1(n1734), .A0N(\gbuff[6][5] ), .A1N(n1736), 
        .Y(n2621) );
  OAI2BB2XL U1003 ( .B0(n1505), .B1(n1734), .A0N(\gbuff[6][6] ), .A1N(n1736), 
        .Y(n2620) );
  OAI2BB2XL U1004 ( .B0(n1503), .B1(n1734), .A0N(\gbuff[6][7] ), .A1N(n1736), 
        .Y(n2619) );
  OAI2BB2XL U1005 ( .B0(n1501), .B1(n1734), .A0N(\gbuff[6][8] ), .A1N(n1736), 
        .Y(n2618) );
  OAI2BB2XL U1006 ( .B0(n1499), .B1(n1734), .A0N(\gbuff[6][9] ), .A1N(n1736), 
        .Y(n2617) );
  OAI2BB2XL U1007 ( .B0(n1497), .B1(n1734), .A0N(\gbuff[6][10] ), .A1N(n1736), 
        .Y(n2616) );
  OAI2BB2XL U1008 ( .B0(n1495), .B1(n1734), .A0N(\gbuff[6][11] ), .A1N(n1736), 
        .Y(n2615) );
  OAI2BB2XL U1009 ( .B0(n1493), .B1(n1734), .A0N(\gbuff[6][12] ), .A1N(n1736), 
        .Y(n2614) );
  OAI2BB2XL U1010 ( .B0(n1491), .B1(n1734), .A0N(\gbuff[6][13] ), .A1N(n1736), 
        .Y(n2613) );
  OAI2BB2XL U1011 ( .B0(n1489), .B1(n1735), .A0N(\gbuff[6][14] ), .A1N(n1736), 
        .Y(n2612) );
  OAI2BB2XL U1012 ( .B0(n1487), .B1(n1734), .A0N(\gbuff[6][15] ), .A1N(n1735), 
        .Y(n2611) );
  OAI2BB2XL U1013 ( .B0(n1485), .B1(n1735), .A0N(\gbuff[6][16] ), .A1N(n1736), 
        .Y(n2610) );
  OAI2BB2XL U1014 ( .B0(n1483), .B1(n1734), .A0N(\gbuff[6][17] ), .A1N(n1735), 
        .Y(n2609) );
  OAI2BB2XL U1015 ( .B0(n1481), .B1(n1735), .A0N(\gbuff[6][18] ), .A1N(n1735), 
        .Y(n2608) );
  OAI2BB2XL U1016 ( .B0(n1479), .B1(n1734), .A0N(\gbuff[6][19] ), .A1N(n1735), 
        .Y(n2607) );
  OAI2BB2XL U1017 ( .B0(n1477), .B1(n1735), .A0N(\gbuff[6][20] ), .A1N(n1735), 
        .Y(n2606) );
  OAI2BB2XL U1018 ( .B0(n1475), .B1(n1734), .A0N(\gbuff[6][21] ), .A1N(n1735), 
        .Y(n2605) );
  OAI2BB2XL U1019 ( .B0(n1473), .B1(n1735), .A0N(\gbuff[6][22] ), .A1N(n1736), 
        .Y(n2604) );
  OAI2BB2XL U1020 ( .B0(n1471), .B1(n1735), .A0N(\gbuff[6][23] ), .A1N(n1735), 
        .Y(n2603) );
  OAI2BB2XL U1021 ( .B0(n1469), .B1(n7), .A0N(\gbuff[6][24] ), .A1N(n1736), 
        .Y(n2602) );
  OAI2BB2XL U1022 ( .B0(n1467), .B1(n1735), .A0N(\gbuff[6][25] ), .A1N(n1736), 
        .Y(n2601) );
  OAI2BB2XL U1023 ( .B0(n1465), .B1(n1735), .A0N(\gbuff[6][26] ), .A1N(n1736), 
        .Y(n2600) );
  OAI2BB2XL U1024 ( .B0(n1463), .B1(n1735), .A0N(\gbuff[6][27] ), .A1N(n1736), 
        .Y(n2599) );
  OAI2BB2XL U1025 ( .B0(n1461), .B1(n1735), .A0N(\gbuff[6][28] ), .A1N(n1736), 
        .Y(n2598) );
  OAI2BB2XL U1026 ( .B0(n1459), .B1(n1735), .A0N(\gbuff[6][29] ), .A1N(n1736), 
        .Y(n2597) );
  OAI2BB2XL U1027 ( .B0(n1457), .B1(n1735), .A0N(\gbuff[6][30] ), .A1N(n1736), 
        .Y(n2596) );
  OAI2BB2XL U1028 ( .B0(n1455), .B1(n1735), .A0N(\gbuff[6][31] ), .A1N(n1734), 
        .Y(n2595) );
  OAI2BB2XL U1029 ( .B0(n1516), .B1(n1731), .A0N(\gbuff[7][0] ), .A1N(n1733), 
        .Y(n2594) );
  OAI2BB2XL U1030 ( .B0(n1514), .B1(n1731), .A0N(\gbuff[7][1] ), .A1N(n8), .Y(
        n2593) );
  OAI2BB2XL U1031 ( .B0(n1512), .B1(n1731), .A0N(\gbuff[7][2] ), .A1N(n1731), 
        .Y(n2592) );
  OAI2BB2XL U1032 ( .B0(n1510), .B1(n1731), .A0N(\gbuff[7][3] ), .A1N(n1733), 
        .Y(n2591) );
  OAI2BB2XL U1033 ( .B0(n1508), .B1(n1731), .A0N(\gbuff[7][4] ), .A1N(n1733), 
        .Y(n2590) );
  OAI2BB2XL U1034 ( .B0(n1506), .B1(n1731), .A0N(\gbuff[7][5] ), .A1N(n1733), 
        .Y(n2589) );
  OAI2BB2XL U1035 ( .B0(n1504), .B1(n1731), .A0N(\gbuff[7][6] ), .A1N(n1733), 
        .Y(n2588) );
  OAI2BB2XL U1036 ( .B0(n1502), .B1(n1731), .A0N(\gbuff[7][7] ), .A1N(n1733), 
        .Y(n2587) );
  OAI2BB2XL U1037 ( .B0(n1500), .B1(n1731), .A0N(\gbuff[7][8] ), .A1N(n1733), 
        .Y(n2586) );
  OAI2BB2XL U1038 ( .B0(n1498), .B1(n1731), .A0N(\gbuff[7][9] ), .A1N(n1733), 
        .Y(n2585) );
  OAI2BB2XL U1039 ( .B0(n1496), .B1(n1731), .A0N(\gbuff[7][10] ), .A1N(n1733), 
        .Y(n2584) );
  OAI2BB2XL U1040 ( .B0(n1494), .B1(n1731), .A0N(\gbuff[7][11] ), .A1N(n1733), 
        .Y(n2583) );
  OAI2BB2XL U1041 ( .B0(n1492), .B1(n1731), .A0N(\gbuff[7][12] ), .A1N(n1733), 
        .Y(n2582) );
  OAI2BB2XL U1042 ( .B0(n1490), .B1(n1731), .A0N(\gbuff[7][13] ), .A1N(n1733), 
        .Y(n2581) );
  OAI2BB2XL U1043 ( .B0(n1488), .B1(n1732), .A0N(\gbuff[7][14] ), .A1N(n1733), 
        .Y(n2580) );
  OAI2BB2XL U1044 ( .B0(n1486), .B1(n1731), .A0N(\gbuff[7][15] ), .A1N(n1732), 
        .Y(n2579) );
  OAI2BB2XL U1045 ( .B0(n1484), .B1(n1732), .A0N(\gbuff[7][16] ), .A1N(n1733), 
        .Y(n2578) );
  OAI2BB2XL U1046 ( .B0(n1482), .B1(n1731), .A0N(\gbuff[7][17] ), .A1N(n1732), 
        .Y(n2577) );
  OAI2BB2XL U1047 ( .B0(n1480), .B1(n1732), .A0N(\gbuff[7][18] ), .A1N(n1732), 
        .Y(n2576) );
  OAI2BB2XL U1048 ( .B0(n1478), .B1(n1731), .A0N(\gbuff[7][19] ), .A1N(n1732), 
        .Y(n2575) );
  OAI2BB2XL U1049 ( .B0(n1476), .B1(n1732), .A0N(\gbuff[7][20] ), .A1N(n1732), 
        .Y(n2574) );
  OAI2BB2XL U1050 ( .B0(n1474), .B1(n1731), .A0N(\gbuff[7][21] ), .A1N(n1732), 
        .Y(n2573) );
  OAI2BB2XL U1051 ( .B0(n1472), .B1(n1732), .A0N(\gbuff[7][22] ), .A1N(n1733), 
        .Y(n2572) );
  OAI2BB2XL U1052 ( .B0(n1470), .B1(n1732), .A0N(\gbuff[7][23] ), .A1N(n1732), 
        .Y(n2571) );
  OAI2BB2XL U1053 ( .B0(n1468), .B1(n8), .A0N(\gbuff[7][24] ), .A1N(n1733), 
        .Y(n2570) );
  OAI2BB2XL U1054 ( .B0(n1466), .B1(n1732), .A0N(\gbuff[7][25] ), .A1N(n1733), 
        .Y(n2569) );
  OAI2BB2XL U1055 ( .B0(n1464), .B1(n1732), .A0N(\gbuff[7][26] ), .A1N(n1733), 
        .Y(n2568) );
  OAI2BB2XL U1056 ( .B0(n1462), .B1(n1732), .A0N(\gbuff[7][27] ), .A1N(n1733), 
        .Y(n2567) );
  OAI2BB2XL U1057 ( .B0(n1460), .B1(n1732), .A0N(\gbuff[7][28] ), .A1N(n1733), 
        .Y(n2566) );
  OAI2BB2XL U1058 ( .B0(n1458), .B1(n1732), .A0N(\gbuff[7][29] ), .A1N(n1733), 
        .Y(n2565) );
  OAI2BB2XL U1059 ( .B0(n1456), .B1(n1732), .A0N(\gbuff[7][30] ), .A1N(n1733), 
        .Y(n2564) );
  OAI2BB2XL U1060 ( .B0(n1454), .B1(n1732), .A0N(\gbuff[7][31] ), .A1N(n1731), 
        .Y(n2563) );
  OAI2BB2XL U1061 ( .B0(n1517), .B1(n1728), .A0N(\gbuff[8][0] ), .A1N(n1730), 
        .Y(n2562) );
  OAI2BB2XL U1062 ( .B0(n1515), .B1(n1728), .A0N(\gbuff[8][1] ), .A1N(n1729), 
        .Y(n2561) );
  OAI2BB2XL U1063 ( .B0(n1513), .B1(n1728), .A0N(\gbuff[8][2] ), .A1N(n1728), 
        .Y(n2560) );
  OAI2BB2XL U1064 ( .B0(n1511), .B1(n1728), .A0N(\gbuff[8][3] ), .A1N(n1730), 
        .Y(n2559) );
  OAI2BB2XL U1065 ( .B0(n1509), .B1(n1728), .A0N(\gbuff[8][4] ), .A1N(n1730), 
        .Y(n2558) );
  OAI2BB2XL U1066 ( .B0(n1507), .B1(n1728), .A0N(\gbuff[8][5] ), .A1N(n1730), 
        .Y(n2557) );
  OAI2BB2XL U1067 ( .B0(n1505), .B1(n1728), .A0N(\gbuff[8][6] ), .A1N(n1730), 
        .Y(n2556) );
  OAI2BB2XL U1068 ( .B0(n1503), .B1(n1728), .A0N(\gbuff[8][7] ), .A1N(n1730), 
        .Y(n2555) );
  OAI2BB2XL U1069 ( .B0(n1501), .B1(n1728), .A0N(\gbuff[8][8] ), .A1N(n1730), 
        .Y(n2554) );
  OAI2BB2XL U1070 ( .B0(n1499), .B1(n1728), .A0N(\gbuff[8][9] ), .A1N(n1730), 
        .Y(n2553) );
  OAI2BB2XL U1071 ( .B0(n1497), .B1(n1728), .A0N(\gbuff[8][10] ), .A1N(n1730), 
        .Y(n2552) );
  OAI2BB2XL U1072 ( .B0(n1495), .B1(n1728), .A0N(\gbuff[8][11] ), .A1N(n1730), 
        .Y(n2551) );
  OAI2BB2XL U1073 ( .B0(n1493), .B1(n1728), .A0N(\gbuff[8][12] ), .A1N(n1730), 
        .Y(n2550) );
  OAI2BB2XL U1074 ( .B0(n1491), .B1(n1728), .A0N(\gbuff[8][13] ), .A1N(n1730), 
        .Y(n2549) );
  OAI2BB2XL U1075 ( .B0(n1489), .B1(n1729), .A0N(\gbuff[8][14] ), .A1N(n1730), 
        .Y(n2548) );
  OAI2BB2XL U1076 ( .B0(n1487), .B1(n1728), .A0N(\gbuff[8][15] ), .A1N(n1729), 
        .Y(n2547) );
  OAI2BB2XL U1077 ( .B0(n1485), .B1(n1729), .A0N(\gbuff[8][16] ), .A1N(n1730), 
        .Y(n2546) );
  OAI2BB2XL U1078 ( .B0(n1483), .B1(n1728), .A0N(\gbuff[8][17] ), .A1N(n1729), 
        .Y(n2545) );
  OAI2BB2XL U1079 ( .B0(n1481), .B1(n1729), .A0N(\gbuff[8][18] ), .A1N(n1729), 
        .Y(n2544) );
  OAI2BB2XL U1080 ( .B0(n1479), .B1(n1728), .A0N(\gbuff[8][19] ), .A1N(n1729), 
        .Y(n2543) );
  OAI2BB2XL U1081 ( .B0(n1477), .B1(n1729), .A0N(\gbuff[8][20] ), .A1N(n1729), 
        .Y(n2542) );
  OAI2BB2XL U1082 ( .B0(n1475), .B1(n1728), .A0N(\gbuff[8][21] ), .A1N(n1729), 
        .Y(n2541) );
  OAI2BB2XL U1083 ( .B0(n1473), .B1(n1729), .A0N(\gbuff[8][22] ), .A1N(n1730), 
        .Y(n2540) );
  OAI2BB2XL U1084 ( .B0(n1471), .B1(n1729), .A0N(\gbuff[8][23] ), .A1N(n1729), 
        .Y(n2539) );
  OAI2BB2XL U1085 ( .B0(n1469), .B1(n1728), .A0N(\gbuff[8][24] ), .A1N(n1730), 
        .Y(n2538) );
  OAI2BB2XL U1086 ( .B0(n1467), .B1(n1729), .A0N(\gbuff[8][25] ), .A1N(n1730), 
        .Y(n2537) );
  OAI2BB2XL U1087 ( .B0(n1465), .B1(n1729), .A0N(\gbuff[8][26] ), .A1N(n1730), 
        .Y(n2536) );
  OAI2BB2XL U1088 ( .B0(n1463), .B1(n1729), .A0N(\gbuff[8][27] ), .A1N(n1730), 
        .Y(n2535) );
  OAI2BB2XL U1089 ( .B0(n1461), .B1(n1729), .A0N(\gbuff[8][28] ), .A1N(n1730), 
        .Y(n2534) );
  OAI2BB2XL U1090 ( .B0(n1459), .B1(n1729), .A0N(\gbuff[8][29] ), .A1N(n1730), 
        .Y(n2533) );
  OAI2BB2XL U1091 ( .B0(n1457), .B1(n1729), .A0N(\gbuff[8][30] ), .A1N(n1730), 
        .Y(n2532) );
  OAI2BB2XL U1092 ( .B0(n1455), .B1(n1729), .A0N(\gbuff[8][31] ), .A1N(n1728), 
        .Y(n2531) );
  OAI2BB2XL U1093 ( .B0(n1517), .B1(n1725), .A0N(\gbuff[9][0] ), .A1N(n1727), 
        .Y(n2530) );
  OAI2BB2XL U1094 ( .B0(n1515), .B1(n1725), .A0N(\gbuff[9][1] ), .A1N(n1726), 
        .Y(n2529) );
  OAI2BB2XL U1095 ( .B0(n1513), .B1(n1725), .A0N(\gbuff[9][2] ), .A1N(n1725), 
        .Y(n2528) );
  OAI2BB2XL U1096 ( .B0(n1511), .B1(n1725), .A0N(\gbuff[9][3] ), .A1N(n1727), 
        .Y(n2527) );
  OAI2BB2XL U1097 ( .B0(n1509), .B1(n1725), .A0N(\gbuff[9][4] ), .A1N(n1727), 
        .Y(n2526) );
  OAI2BB2XL U1098 ( .B0(n1507), .B1(n1725), .A0N(\gbuff[9][5] ), .A1N(n1727), 
        .Y(n2525) );
  OAI2BB2XL U1099 ( .B0(n1505), .B1(n1725), .A0N(\gbuff[9][6] ), .A1N(n1727), 
        .Y(n2524) );
  OAI2BB2XL U1100 ( .B0(n1503), .B1(n1725), .A0N(\gbuff[9][7] ), .A1N(n1727), 
        .Y(n2523) );
  OAI2BB2XL U1101 ( .B0(n1501), .B1(n1725), .A0N(\gbuff[9][8] ), .A1N(n1727), 
        .Y(n2522) );
  OAI2BB2XL U1102 ( .B0(n1499), .B1(n1725), .A0N(\gbuff[9][9] ), .A1N(n1727), 
        .Y(n2521) );
  OAI2BB2XL U1103 ( .B0(n1497), .B1(n1725), .A0N(\gbuff[9][10] ), .A1N(n1727), 
        .Y(n2520) );
  OAI2BB2XL U1104 ( .B0(n1495), .B1(n1725), .A0N(\gbuff[9][11] ), .A1N(n1727), 
        .Y(n2519) );
  OAI2BB2XL U1105 ( .B0(n1493), .B1(n1725), .A0N(\gbuff[9][12] ), .A1N(n1727), 
        .Y(n2518) );
  OAI2BB2XL U1106 ( .B0(n1491), .B1(n1725), .A0N(\gbuff[9][13] ), .A1N(n1727), 
        .Y(n2517) );
  OAI2BB2XL U1107 ( .B0(n1489), .B1(n1726), .A0N(\gbuff[9][14] ), .A1N(n1727), 
        .Y(n2516) );
  OAI2BB2XL U1108 ( .B0(n1487), .B1(n1725), .A0N(\gbuff[9][15] ), .A1N(n1726), 
        .Y(n2515) );
  OAI2BB2XL U1109 ( .B0(n1485), .B1(n1726), .A0N(\gbuff[9][16] ), .A1N(n1727), 
        .Y(n2514) );
  OAI2BB2XL U1110 ( .B0(n1483), .B1(n1725), .A0N(\gbuff[9][17] ), .A1N(n1726), 
        .Y(n2513) );
  OAI2BB2XL U1111 ( .B0(n1481), .B1(n1726), .A0N(\gbuff[9][18] ), .A1N(n1726), 
        .Y(n2512) );
  OAI2BB2XL U1112 ( .B0(n1479), .B1(n1725), .A0N(\gbuff[9][19] ), .A1N(n1726), 
        .Y(n2511) );
  OAI2BB2XL U1113 ( .B0(n1477), .B1(n1726), .A0N(\gbuff[9][20] ), .A1N(n1726), 
        .Y(n2510) );
  OAI2BB2XL U1114 ( .B0(n1475), .B1(n1725), .A0N(\gbuff[9][21] ), .A1N(n1726), 
        .Y(n2509) );
  OAI2BB2XL U1115 ( .B0(n1473), .B1(n1726), .A0N(\gbuff[9][22] ), .A1N(n1727), 
        .Y(n2508) );
  OAI2BB2XL U1116 ( .B0(n1471), .B1(n1726), .A0N(\gbuff[9][23] ), .A1N(n1726), 
        .Y(n2507) );
  OAI2BB2XL U1117 ( .B0(n1469), .B1(n1725), .A0N(\gbuff[9][24] ), .A1N(n1727), 
        .Y(n2506) );
  OAI2BB2XL U1118 ( .B0(n1467), .B1(n1726), .A0N(\gbuff[9][25] ), .A1N(n1727), 
        .Y(n2505) );
  OAI2BB2XL U1119 ( .B0(n1465), .B1(n1726), .A0N(\gbuff[9][26] ), .A1N(n1727), 
        .Y(n2504) );
  OAI2BB2XL U1120 ( .B0(n1463), .B1(n1726), .A0N(\gbuff[9][27] ), .A1N(n1727), 
        .Y(n2503) );
  OAI2BB2XL U1121 ( .B0(n1461), .B1(n1726), .A0N(\gbuff[9][28] ), .A1N(n1727), 
        .Y(n2502) );
  OAI2BB2XL U1122 ( .B0(n1459), .B1(n1726), .A0N(\gbuff[9][29] ), .A1N(n1727), 
        .Y(n2501) );
  OAI2BB2XL U1123 ( .B0(n1457), .B1(n1726), .A0N(\gbuff[9][30] ), .A1N(n1727), 
        .Y(n2500) );
  OAI2BB2XL U1124 ( .B0(n1455), .B1(n1726), .A0N(\gbuff[9][31] ), .A1N(n1725), 
        .Y(n2499) );
  OAI2BB2XL U1125 ( .B0(n1517), .B1(n1722), .A0N(\gbuff[10][0] ), .A1N(n1724), 
        .Y(n2498) );
  OAI2BB2XL U1126 ( .B0(n1515), .B1(n1722), .A0N(\gbuff[10][1] ), .A1N(n1723), 
        .Y(n2497) );
  OAI2BB2XL U1127 ( .B0(n1513), .B1(n1722), .A0N(\gbuff[10][2] ), .A1N(n1722), 
        .Y(n2496) );
  OAI2BB2XL U1128 ( .B0(n1511), .B1(n1722), .A0N(\gbuff[10][3] ), .A1N(n1724), 
        .Y(n2495) );
  OAI2BB2XL U1129 ( .B0(n1509), .B1(n1722), .A0N(\gbuff[10][4] ), .A1N(n1724), 
        .Y(n2494) );
  OAI2BB2XL U1130 ( .B0(n1507), .B1(n1722), .A0N(\gbuff[10][5] ), .A1N(n1724), 
        .Y(n2493) );
  OAI2BB2XL U1131 ( .B0(n1505), .B1(n1722), .A0N(\gbuff[10][6] ), .A1N(n1724), 
        .Y(n2492) );
  OAI2BB2XL U1132 ( .B0(n1503), .B1(n1722), .A0N(\gbuff[10][7] ), .A1N(n1724), 
        .Y(n2491) );
  OAI2BB2XL U1133 ( .B0(n1501), .B1(n1722), .A0N(\gbuff[10][8] ), .A1N(n1724), 
        .Y(n2490) );
  OAI2BB2XL U1134 ( .B0(n1499), .B1(n1722), .A0N(\gbuff[10][9] ), .A1N(n1724), 
        .Y(n2489) );
  OAI2BB2XL U1135 ( .B0(n1497), .B1(n1722), .A0N(\gbuff[10][10] ), .A1N(n1724), 
        .Y(n2488) );
  OAI2BB2XL U1136 ( .B0(n1495), .B1(n1722), .A0N(\gbuff[10][11] ), .A1N(n1724), 
        .Y(n2487) );
  OAI2BB2XL U1137 ( .B0(n1493), .B1(n1722), .A0N(\gbuff[10][12] ), .A1N(n1724), 
        .Y(n2486) );
  OAI2BB2XL U1138 ( .B0(n1491), .B1(n1722), .A0N(\gbuff[10][13] ), .A1N(n1724), 
        .Y(n2485) );
  OAI2BB2XL U1139 ( .B0(n1489), .B1(n1723), .A0N(\gbuff[10][14] ), .A1N(n1724), 
        .Y(n2484) );
  OAI2BB2XL U1140 ( .B0(n1487), .B1(n1722), .A0N(\gbuff[10][15] ), .A1N(n1723), 
        .Y(n2483) );
  OAI2BB2XL U1141 ( .B0(n1485), .B1(n1723), .A0N(\gbuff[10][16] ), .A1N(n1724), 
        .Y(n2482) );
  OAI2BB2XL U1142 ( .B0(n1483), .B1(n1722), .A0N(\gbuff[10][17] ), .A1N(n1723), 
        .Y(n2481) );
  OAI2BB2XL U1143 ( .B0(n1481), .B1(n1723), .A0N(\gbuff[10][18] ), .A1N(n1723), 
        .Y(n2480) );
  OAI2BB2XL U1144 ( .B0(n1479), .B1(n1722), .A0N(\gbuff[10][19] ), .A1N(n1723), 
        .Y(n2479) );
  OAI2BB2XL U1145 ( .B0(n1477), .B1(n1723), .A0N(\gbuff[10][20] ), .A1N(n1723), 
        .Y(n2478) );
  OAI2BB2XL U1146 ( .B0(n1475), .B1(n1722), .A0N(\gbuff[10][21] ), .A1N(n1723), 
        .Y(n2477) );
  OAI2BB2XL U1147 ( .B0(n1473), .B1(n1723), .A0N(\gbuff[10][22] ), .A1N(n1724), 
        .Y(n2476) );
  OAI2BB2XL U1148 ( .B0(n1471), .B1(n1723), .A0N(\gbuff[10][23] ), .A1N(n1723), 
        .Y(n2475) );
  OAI2BB2XL U1149 ( .B0(n1469), .B1(n1722), .A0N(\gbuff[10][24] ), .A1N(n1724), 
        .Y(n2474) );
  OAI2BB2XL U1150 ( .B0(n1467), .B1(n1723), .A0N(\gbuff[10][25] ), .A1N(n1724), 
        .Y(n2473) );
  OAI2BB2XL U1151 ( .B0(n1465), .B1(n1723), .A0N(\gbuff[10][26] ), .A1N(n1724), 
        .Y(n2472) );
  OAI2BB2XL U1152 ( .B0(n1463), .B1(n1723), .A0N(\gbuff[10][27] ), .A1N(n1724), 
        .Y(n2471) );
  OAI2BB2XL U1153 ( .B0(n1461), .B1(n1723), .A0N(\gbuff[10][28] ), .A1N(n1724), 
        .Y(n2470) );
  OAI2BB2XL U1154 ( .B0(n1459), .B1(n1723), .A0N(\gbuff[10][29] ), .A1N(n1724), 
        .Y(n2469) );
  OAI2BB2XL U1155 ( .B0(n1457), .B1(n1723), .A0N(\gbuff[10][30] ), .A1N(n1724), 
        .Y(n2468) );
  OAI2BB2XL U1156 ( .B0(n1455), .B1(n1723), .A0N(\gbuff[10][31] ), .A1N(n1722), 
        .Y(n2467) );
  OAI2BB2XL U1157 ( .B0(n1517), .B1(n1719), .A0N(\gbuff[11][0] ), .A1N(n1721), 
        .Y(n2466) );
  OAI2BB2XL U1158 ( .B0(n1515), .B1(n1719), .A0N(\gbuff[11][1] ), .A1N(n1720), 
        .Y(n2465) );
  OAI2BB2XL U1159 ( .B0(n1513), .B1(n1719), .A0N(\gbuff[11][2] ), .A1N(n1719), 
        .Y(n2464) );
  OAI2BB2XL U1160 ( .B0(n1511), .B1(n1719), .A0N(\gbuff[11][3] ), .A1N(n1721), 
        .Y(n2463) );
  OAI2BB2XL U1161 ( .B0(n1509), .B1(n1719), .A0N(\gbuff[11][4] ), .A1N(n1721), 
        .Y(n2462) );
  OAI2BB2XL U1162 ( .B0(n1507), .B1(n1719), .A0N(\gbuff[11][5] ), .A1N(n1721), 
        .Y(n2461) );
  OAI2BB2XL U1163 ( .B0(n1505), .B1(n1719), .A0N(\gbuff[11][6] ), .A1N(n1721), 
        .Y(n2460) );
  OAI2BB2XL U1164 ( .B0(n1503), .B1(n1719), .A0N(\gbuff[11][7] ), .A1N(n1721), 
        .Y(n2459) );
  OAI2BB2XL U1165 ( .B0(n1501), .B1(n1719), .A0N(\gbuff[11][8] ), .A1N(n1721), 
        .Y(n2458) );
  OAI2BB2XL U1166 ( .B0(n1499), .B1(n1719), .A0N(\gbuff[11][9] ), .A1N(n1721), 
        .Y(n2457) );
  OAI2BB2XL U1167 ( .B0(n1497), .B1(n1719), .A0N(\gbuff[11][10] ), .A1N(n1721), 
        .Y(n2456) );
  OAI2BB2XL U1168 ( .B0(n1495), .B1(n1719), .A0N(\gbuff[11][11] ), .A1N(n1721), 
        .Y(n2455) );
  OAI2BB2XL U1169 ( .B0(n1493), .B1(n1719), .A0N(\gbuff[11][12] ), .A1N(n1721), 
        .Y(n2454) );
  OAI2BB2XL U1170 ( .B0(n1491), .B1(n1719), .A0N(\gbuff[11][13] ), .A1N(n1721), 
        .Y(n2453) );
  OAI2BB2XL U1171 ( .B0(n1489), .B1(n1720), .A0N(\gbuff[11][14] ), .A1N(n1721), 
        .Y(n2452) );
  OAI2BB2XL U1172 ( .B0(n1487), .B1(n1719), .A0N(\gbuff[11][15] ), .A1N(n1720), 
        .Y(n2451) );
  OAI2BB2XL U1173 ( .B0(n1485), .B1(n1720), .A0N(\gbuff[11][16] ), .A1N(n1721), 
        .Y(n2450) );
  OAI2BB2XL U1174 ( .B0(n1483), .B1(n1719), .A0N(\gbuff[11][17] ), .A1N(n1720), 
        .Y(n2449) );
  OAI2BB2XL U1175 ( .B0(n1481), .B1(n1720), .A0N(\gbuff[11][18] ), .A1N(n1720), 
        .Y(n2448) );
  OAI2BB2XL U1176 ( .B0(n1479), .B1(n1719), .A0N(\gbuff[11][19] ), .A1N(n1720), 
        .Y(n2447) );
  OAI2BB2XL U1177 ( .B0(n1477), .B1(n1720), .A0N(\gbuff[11][20] ), .A1N(n1720), 
        .Y(n2446) );
  OAI2BB2XL U1178 ( .B0(n1475), .B1(n1719), .A0N(\gbuff[11][21] ), .A1N(n1720), 
        .Y(n2445) );
  OAI2BB2XL U1179 ( .B0(n1473), .B1(n1720), .A0N(\gbuff[11][22] ), .A1N(n1721), 
        .Y(n2444) );
  OAI2BB2XL U1180 ( .B0(n1471), .B1(n1720), .A0N(\gbuff[11][23] ), .A1N(n1720), 
        .Y(n2443) );
  OAI2BB2XL U1181 ( .B0(n1469), .B1(n1719), .A0N(\gbuff[11][24] ), .A1N(n1721), 
        .Y(n2442) );
  OAI2BB2XL U1182 ( .B0(n1467), .B1(n1720), .A0N(\gbuff[11][25] ), .A1N(n1721), 
        .Y(n2441) );
  OAI2BB2XL U1183 ( .B0(n1465), .B1(n1720), .A0N(\gbuff[11][26] ), .A1N(n1721), 
        .Y(n2440) );
  OAI2BB2XL U1184 ( .B0(n1463), .B1(n1720), .A0N(\gbuff[11][27] ), .A1N(n1721), 
        .Y(n2439) );
  OAI2BB2XL U1185 ( .B0(n1461), .B1(n1720), .A0N(\gbuff[11][28] ), .A1N(n1721), 
        .Y(n2438) );
  OAI2BB2XL U1186 ( .B0(n1459), .B1(n1720), .A0N(\gbuff[11][29] ), .A1N(n1721), 
        .Y(n2437) );
  OAI2BB2XL U1187 ( .B0(n1457), .B1(n1720), .A0N(\gbuff[11][30] ), .A1N(n1721), 
        .Y(n2436) );
  OAI2BB2XL U1188 ( .B0(n1455), .B1(n1720), .A0N(\gbuff[11][31] ), .A1N(n1719), 
        .Y(n2435) );
  OAI2BB2XL U1189 ( .B0(n1517), .B1(n1717), .A0N(\gbuff[12][0] ), .A1N(n1717), 
        .Y(n2434) );
  OAI2BB2XL U1190 ( .B0(n1515), .B1(n1716), .A0N(\gbuff[12][1] ), .A1N(n1716), 
        .Y(n2433) );
  OAI2BB2XL U1191 ( .B0(n1513), .B1(n1716), .A0N(\gbuff[12][2] ), .A1N(n1717), 
        .Y(n2432) );
  OAI2BB2XL U1192 ( .B0(n1511), .B1(n1716), .A0N(\gbuff[12][3] ), .A1N(n1718), 
        .Y(n2431) );
  OAI2BB2XL U1193 ( .B0(n1509), .B1(n1716), .A0N(\gbuff[12][4] ), .A1N(n1716), 
        .Y(n2430) );
  OAI2BB2XL U1194 ( .B0(n1507), .B1(n1716), .A0N(\gbuff[12][5] ), .A1N(n1718), 
        .Y(n2429) );
  OAI2BB2XL U1195 ( .B0(n1505), .B1(n1716), .A0N(\gbuff[12][6] ), .A1N(n1718), 
        .Y(n2428) );
  OAI2BB2XL U1196 ( .B0(n1503), .B1(n1716), .A0N(\gbuff[12][7] ), .A1N(n1718), 
        .Y(n2427) );
  OAI2BB2XL U1197 ( .B0(n1501), .B1(n1716), .A0N(\gbuff[12][8] ), .A1N(n1718), 
        .Y(n2426) );
  OAI2BB2XL U1198 ( .B0(n1499), .B1(n1716), .A0N(\gbuff[12][9] ), .A1N(n1718), 
        .Y(n2425) );
  OAI2BB2XL U1199 ( .B0(n1497), .B1(n1716), .A0N(\gbuff[12][10] ), .A1N(n1718), 
        .Y(n2424) );
  OAI2BB2XL U1200 ( .B0(n1495), .B1(n1716), .A0N(\gbuff[12][11] ), .A1N(n1718), 
        .Y(n2423) );
  OAI2BB2XL U1201 ( .B0(n1493), .B1(n1716), .A0N(\gbuff[12][12] ), .A1N(n1718), 
        .Y(n2422) );
  OAI2BB2XL U1202 ( .B0(n1491), .B1(n1717), .A0N(\gbuff[12][13] ), .A1N(n1718), 
        .Y(n2421) );
  OAI2BB2XL U1203 ( .B0(n1489), .B1(n1717), .A0N(\gbuff[12][14] ), .A1N(n1718), 
        .Y(n2420) );
  OAI2BB2XL U1204 ( .B0(n1487), .B1(n1717), .A0N(\gbuff[12][15] ), .A1N(n1717), 
        .Y(n2419) );
  OAI2BB2XL U1205 ( .B0(n1485), .B1(n1717), .A0N(\gbuff[12][16] ), .A1N(n1718), 
        .Y(n2418) );
  OAI2BB2XL U1206 ( .B0(n1483), .B1(n1717), .A0N(\gbuff[12][17] ), .A1N(n1716), 
        .Y(n2417) );
  OAI2BB2XL U1207 ( .B0(n1481), .B1(n1717), .A0N(\gbuff[12][18] ), .A1N(n1718), 
        .Y(n2416) );
  OAI2BB2XL U1208 ( .B0(n1479), .B1(n1717), .A0N(\gbuff[12][19] ), .A1N(n1717), 
        .Y(n2415) );
  OAI2BB2XL U1209 ( .B0(n1477), .B1(n1717), .A0N(\gbuff[12][20] ), .A1N(n1716), 
        .Y(n2414) );
  OAI2BB2XL U1210 ( .B0(n1475), .B1(n1717), .A0N(\gbuff[12][21] ), .A1N(n1718), 
        .Y(n2413) );
  OAI2BB2XL U1211 ( .B0(n1473), .B1(n1717), .A0N(\gbuff[12][22] ), .A1N(n1718), 
        .Y(n2412) );
  OAI2BB2XL U1212 ( .B0(n1471), .B1(n1717), .A0N(\gbuff[12][23] ), .A1N(n1718), 
        .Y(n2411) );
  OAI2BB2XL U1213 ( .B0(n1469), .B1(n1717), .A0N(\gbuff[12][24] ), .A1N(n1718), 
        .Y(n2410) );
  OAI2BB2XL U1214 ( .B0(n1467), .B1(n1716), .A0N(\gbuff[12][25] ), .A1N(n1718), 
        .Y(n2409) );
  OAI2BB2XL U1215 ( .B0(n1465), .B1(n1717), .A0N(\gbuff[12][26] ), .A1N(n1718), 
        .Y(n2408) );
  OAI2BB2XL U1216 ( .B0(n1463), .B1(n1716), .A0N(\gbuff[12][27] ), .A1N(n1718), 
        .Y(n2407) );
  OAI2BB2XL U1217 ( .B0(n1461), .B1(n1717), .A0N(\gbuff[12][28] ), .A1N(n1718), 
        .Y(n2406) );
  OAI2BB2XL U1218 ( .B0(n1459), .B1(n1716), .A0N(\gbuff[12][29] ), .A1N(n1718), 
        .Y(n2405) );
  OAI2BB2XL U1219 ( .B0(n1457), .B1(n1717), .A0N(\gbuff[12][30] ), .A1N(n1717), 
        .Y(n2404) );
  OAI2BB2XL U1220 ( .B0(n1455), .B1(n1716), .A0N(\gbuff[12][31] ), .A1N(n1716), 
        .Y(n2403) );
  OAI2BB2XL U1221 ( .B0(n1517), .B1(n1713), .A0N(\gbuff[13][0] ), .A1N(n1715), 
        .Y(n2402) );
  OAI2BB2XL U1222 ( .B0(n1515), .B1(n1713), .A0N(\gbuff[13][1] ), .A1N(n14), 
        .Y(n2401) );
  OAI2BB2XL U1223 ( .B0(n1513), .B1(n1713), .A0N(\gbuff[13][2] ), .A1N(n1713), 
        .Y(n2400) );
  OAI2BB2XL U1224 ( .B0(n1511), .B1(n1713), .A0N(\gbuff[13][3] ), .A1N(n1715), 
        .Y(n2399) );
  OAI2BB2XL U1225 ( .B0(n1509), .B1(n1713), .A0N(\gbuff[13][4] ), .A1N(n1715), 
        .Y(n2398) );
  OAI2BB2XL U1226 ( .B0(n1507), .B1(n1713), .A0N(\gbuff[13][5] ), .A1N(n1715), 
        .Y(n2397) );
  OAI2BB2XL U1227 ( .B0(n1505), .B1(n1713), .A0N(\gbuff[13][6] ), .A1N(n1715), 
        .Y(n2396) );
  OAI2BB2XL U1228 ( .B0(n1503), .B1(n1713), .A0N(\gbuff[13][7] ), .A1N(n1715), 
        .Y(n2395) );
  OAI2BB2XL U1229 ( .B0(n1501), .B1(n1713), .A0N(\gbuff[13][8] ), .A1N(n1715), 
        .Y(n2394) );
  OAI2BB2XL U1230 ( .B0(n1499), .B1(n1713), .A0N(\gbuff[13][9] ), .A1N(n1715), 
        .Y(n2393) );
  OAI2BB2XL U1231 ( .B0(n1497), .B1(n1713), .A0N(\gbuff[13][10] ), .A1N(n1715), 
        .Y(n2392) );
  OAI2BB2XL U1232 ( .B0(n1495), .B1(n1713), .A0N(\gbuff[13][11] ), .A1N(n1715), 
        .Y(n2391) );
  OAI2BB2XL U1233 ( .B0(n1493), .B1(n1713), .A0N(\gbuff[13][12] ), .A1N(n1715), 
        .Y(n2390) );
  OAI2BB2XL U1234 ( .B0(n1491), .B1(n1713), .A0N(\gbuff[13][13] ), .A1N(n1715), 
        .Y(n2389) );
  OAI2BB2XL U1235 ( .B0(n1489), .B1(n1714), .A0N(\gbuff[13][14] ), .A1N(n1715), 
        .Y(n2388) );
  OAI2BB2XL U1236 ( .B0(n1487), .B1(n1713), .A0N(\gbuff[13][15] ), .A1N(n1714), 
        .Y(n2387) );
  OAI2BB2XL U1237 ( .B0(n1485), .B1(n1714), .A0N(\gbuff[13][16] ), .A1N(n1715), 
        .Y(n2386) );
  OAI2BB2XL U1238 ( .B0(n1483), .B1(n1713), .A0N(\gbuff[13][17] ), .A1N(n1714), 
        .Y(n2385) );
  OAI2BB2XL U1239 ( .B0(n1481), .B1(n1714), .A0N(\gbuff[13][18] ), .A1N(n1714), 
        .Y(n2384) );
  OAI2BB2XL U1240 ( .B0(n1479), .B1(n1713), .A0N(\gbuff[13][19] ), .A1N(n1714), 
        .Y(n2383) );
  OAI2BB2XL U1241 ( .B0(n1477), .B1(n1714), .A0N(\gbuff[13][20] ), .A1N(n1714), 
        .Y(n2382) );
  OAI2BB2XL U1242 ( .B0(n1475), .B1(n1713), .A0N(\gbuff[13][21] ), .A1N(n1714), 
        .Y(n2381) );
  OAI2BB2XL U1243 ( .B0(n1473), .B1(n1714), .A0N(\gbuff[13][22] ), .A1N(n1715), 
        .Y(n2380) );
  OAI2BB2XL U1244 ( .B0(n1471), .B1(n1714), .A0N(\gbuff[13][23] ), .A1N(n1714), 
        .Y(n2379) );
  OAI2BB2XL U1245 ( .B0(n1469), .B1(n14), .A0N(\gbuff[13][24] ), .A1N(n1715), 
        .Y(n2378) );
  OAI2BB2XL U1246 ( .B0(n1467), .B1(n1714), .A0N(\gbuff[13][25] ), .A1N(n1715), 
        .Y(n2377) );
  OAI2BB2XL U1247 ( .B0(n1465), .B1(n1714), .A0N(\gbuff[13][26] ), .A1N(n1715), 
        .Y(n2376) );
  OAI2BB2XL U1248 ( .B0(n1463), .B1(n1714), .A0N(\gbuff[13][27] ), .A1N(n1715), 
        .Y(n2375) );
  OAI2BB2XL U1249 ( .B0(n1461), .B1(n1714), .A0N(\gbuff[13][28] ), .A1N(n1715), 
        .Y(n2374) );
  OAI2BB2XL U1250 ( .B0(n1459), .B1(n1714), .A0N(\gbuff[13][29] ), .A1N(n1715), 
        .Y(n2373) );
  OAI2BB2XL U1251 ( .B0(n1457), .B1(n1714), .A0N(\gbuff[13][30] ), .A1N(n1715), 
        .Y(n2372) );
  OAI2BB2XL U1252 ( .B0(n1455), .B1(n1714), .A0N(\gbuff[13][31] ), .A1N(n1713), 
        .Y(n2371) );
  OAI2BB2XL U1253 ( .B0(n1517), .B1(n1710), .A0N(\gbuff[14][0] ), .A1N(n1712), 
        .Y(n2370) );
  OAI2BB2XL U1254 ( .B0(n1515), .B1(n1710), .A0N(\gbuff[14][1] ), .A1N(n15), 
        .Y(n2369) );
  OAI2BB2XL U1255 ( .B0(n1513), .B1(n1710), .A0N(\gbuff[14][2] ), .A1N(n1710), 
        .Y(n2368) );
  OAI2BB2XL U1256 ( .B0(n1511), .B1(n1710), .A0N(\gbuff[14][3] ), .A1N(n1712), 
        .Y(n2367) );
  OAI2BB2XL U1257 ( .B0(n1509), .B1(n1710), .A0N(\gbuff[14][4] ), .A1N(n1712), 
        .Y(n2366) );
  OAI2BB2XL U1258 ( .B0(n1507), .B1(n1710), .A0N(\gbuff[14][5] ), .A1N(n1712), 
        .Y(n2365) );
  OAI2BB2XL U1259 ( .B0(n1505), .B1(n1710), .A0N(\gbuff[14][6] ), .A1N(n1712), 
        .Y(n2364) );
  OAI2BB2XL U1260 ( .B0(n1503), .B1(n1710), .A0N(\gbuff[14][7] ), .A1N(n1712), 
        .Y(n2363) );
  OAI2BB2XL U1261 ( .B0(n1501), .B1(n1710), .A0N(\gbuff[14][8] ), .A1N(n1712), 
        .Y(n2362) );
  OAI2BB2XL U1262 ( .B0(n1499), .B1(n1710), .A0N(\gbuff[14][9] ), .A1N(n1712), 
        .Y(n2361) );
  OAI2BB2XL U1263 ( .B0(n1497), .B1(n1710), .A0N(\gbuff[14][10] ), .A1N(n1712), 
        .Y(n2360) );
  OAI2BB2XL U1264 ( .B0(n1495), .B1(n1710), .A0N(\gbuff[14][11] ), .A1N(n1712), 
        .Y(n2359) );
  OAI2BB2XL U1265 ( .B0(n1493), .B1(n1710), .A0N(\gbuff[14][12] ), .A1N(n1712), 
        .Y(n2358) );
  OAI2BB2XL U1266 ( .B0(n1491), .B1(n1710), .A0N(\gbuff[14][13] ), .A1N(n1712), 
        .Y(n2357) );
  OAI2BB2XL U1267 ( .B0(n1489), .B1(n1711), .A0N(\gbuff[14][14] ), .A1N(n1712), 
        .Y(n2356) );
  OAI2BB2XL U1268 ( .B0(n1487), .B1(n1710), .A0N(\gbuff[14][15] ), .A1N(n1711), 
        .Y(n2355) );
  OAI2BB2XL U1269 ( .B0(n1485), .B1(n1711), .A0N(\gbuff[14][16] ), .A1N(n1712), 
        .Y(n2354) );
  OAI2BB2XL U1270 ( .B0(n1483), .B1(n1710), .A0N(\gbuff[14][17] ), .A1N(n1711), 
        .Y(n2353) );
  OAI2BB2XL U1271 ( .B0(n1481), .B1(n1711), .A0N(\gbuff[14][18] ), .A1N(n1711), 
        .Y(n2352) );
  OAI2BB2XL U1272 ( .B0(n1479), .B1(n1710), .A0N(\gbuff[14][19] ), .A1N(n1711), 
        .Y(n2351) );
  OAI2BB2XL U1273 ( .B0(n1477), .B1(n1711), .A0N(\gbuff[14][20] ), .A1N(n1711), 
        .Y(n2350) );
  OAI2BB2XL U1274 ( .B0(n1475), .B1(n1710), .A0N(\gbuff[14][21] ), .A1N(n1711), 
        .Y(n2349) );
  OAI2BB2XL U1275 ( .B0(n1473), .B1(n1711), .A0N(\gbuff[14][22] ), .A1N(n1712), 
        .Y(n2348) );
  OAI2BB2XL U1276 ( .B0(n1471), .B1(n1711), .A0N(\gbuff[14][23] ), .A1N(n1711), 
        .Y(n2347) );
  OAI2BB2XL U1277 ( .B0(n1469), .B1(n15), .A0N(\gbuff[14][24] ), .A1N(n1712), 
        .Y(n2346) );
  OAI2BB2XL U1278 ( .B0(n1467), .B1(n1711), .A0N(\gbuff[14][25] ), .A1N(n1712), 
        .Y(n2345) );
  OAI2BB2XL U1279 ( .B0(n1465), .B1(n1711), .A0N(\gbuff[14][26] ), .A1N(n1712), 
        .Y(n2344) );
  OAI2BB2XL U1280 ( .B0(n1463), .B1(n1711), .A0N(\gbuff[14][27] ), .A1N(n1712), 
        .Y(n2343) );
  OAI2BB2XL U1281 ( .B0(n1461), .B1(n1711), .A0N(\gbuff[14][28] ), .A1N(n1712), 
        .Y(n2342) );
  OAI2BB2XL U1282 ( .B0(n1459), .B1(n1711), .A0N(\gbuff[14][29] ), .A1N(n1712), 
        .Y(n2341) );
  OAI2BB2XL U1283 ( .B0(n1457), .B1(n1711), .A0N(\gbuff[14][30] ), .A1N(n1712), 
        .Y(n2340) );
  OAI2BB2XL U1284 ( .B0(n1455), .B1(n1711), .A0N(\gbuff[14][31] ), .A1N(n1710), 
        .Y(n2339) );
  OAI2BB2XL U1285 ( .B0(n1517), .B1(n1707), .A0N(\gbuff[15][0] ), .A1N(n1709), 
        .Y(n2338) );
  OAI2BB2XL U1286 ( .B0(n1515), .B1(n1707), .A0N(\gbuff[15][1] ), .A1N(n16), 
        .Y(n2337) );
  OAI2BB2XL U1287 ( .B0(n1513), .B1(n1707), .A0N(\gbuff[15][2] ), .A1N(n1707), 
        .Y(n2336) );
  OAI2BB2XL U1288 ( .B0(n1511), .B1(n1707), .A0N(\gbuff[15][3] ), .A1N(n1709), 
        .Y(n2335) );
  OAI2BB2XL U1289 ( .B0(n1509), .B1(n1707), .A0N(\gbuff[15][4] ), .A1N(n1709), 
        .Y(n2334) );
  OAI2BB2XL U1290 ( .B0(n1507), .B1(n1707), .A0N(\gbuff[15][5] ), .A1N(n1709), 
        .Y(n2333) );
  OAI2BB2XL U1291 ( .B0(n1505), .B1(n1707), .A0N(\gbuff[15][6] ), .A1N(n1709), 
        .Y(n2332) );
  OAI2BB2XL U1292 ( .B0(n1503), .B1(n1707), .A0N(\gbuff[15][7] ), .A1N(n1709), 
        .Y(n2331) );
  OAI2BB2XL U1293 ( .B0(n1501), .B1(n1707), .A0N(\gbuff[15][8] ), .A1N(n1709), 
        .Y(n2330) );
  OAI2BB2XL U1294 ( .B0(n1499), .B1(n1707), .A0N(\gbuff[15][9] ), .A1N(n1709), 
        .Y(n2329) );
  OAI2BB2XL U1295 ( .B0(n1497), .B1(n1707), .A0N(\gbuff[15][10] ), .A1N(n1709), 
        .Y(n2328) );
  OAI2BB2XL U1296 ( .B0(n1495), .B1(n1707), .A0N(\gbuff[15][11] ), .A1N(n1709), 
        .Y(n2327) );
  OAI2BB2XL U1297 ( .B0(n1493), .B1(n1707), .A0N(\gbuff[15][12] ), .A1N(n1709), 
        .Y(n2326) );
  OAI2BB2XL U1298 ( .B0(n1491), .B1(n1707), .A0N(\gbuff[15][13] ), .A1N(n1709), 
        .Y(n2325) );
  OAI2BB2XL U1299 ( .B0(n1489), .B1(n1708), .A0N(\gbuff[15][14] ), .A1N(n1709), 
        .Y(n2324) );
  OAI2BB2XL U1300 ( .B0(n1487), .B1(n1707), .A0N(\gbuff[15][15] ), .A1N(n1708), 
        .Y(n2323) );
  OAI2BB2XL U1301 ( .B0(n1485), .B1(n1708), .A0N(\gbuff[15][16] ), .A1N(n1709), 
        .Y(n2322) );
  OAI2BB2XL U1302 ( .B0(n1483), .B1(n1707), .A0N(\gbuff[15][17] ), .A1N(n1708), 
        .Y(n2321) );
  OAI2BB2XL U1303 ( .B0(n1481), .B1(n1708), .A0N(\gbuff[15][18] ), .A1N(n1708), 
        .Y(n2320) );
  OAI2BB2XL U1304 ( .B0(n1479), .B1(n1707), .A0N(\gbuff[15][19] ), .A1N(n1708), 
        .Y(n2319) );
  OAI2BB2XL U1305 ( .B0(n1477), .B1(n1708), .A0N(\gbuff[15][20] ), .A1N(n1708), 
        .Y(n2318) );
  OAI2BB2XL U1306 ( .B0(n1475), .B1(n1707), .A0N(\gbuff[15][21] ), .A1N(n1708), 
        .Y(n2317) );
  OAI2BB2XL U1307 ( .B0(n1473), .B1(n1708), .A0N(\gbuff[15][22] ), .A1N(n1709), 
        .Y(n2316) );
  OAI2BB2XL U1308 ( .B0(n1471), .B1(n1708), .A0N(\gbuff[15][23] ), .A1N(n1708), 
        .Y(n2315) );
  OAI2BB2XL U1309 ( .B0(n1469), .B1(n16), .A0N(\gbuff[15][24] ), .A1N(n1709), 
        .Y(n2314) );
  OAI2BB2XL U1310 ( .B0(n1467), .B1(n1708), .A0N(\gbuff[15][25] ), .A1N(n1709), 
        .Y(n2313) );
  OAI2BB2XL U1311 ( .B0(n1465), .B1(n1708), .A0N(\gbuff[15][26] ), .A1N(n1709), 
        .Y(n2312) );
  OAI2BB2XL U1312 ( .B0(n1463), .B1(n1708), .A0N(\gbuff[15][27] ), .A1N(n1709), 
        .Y(n2311) );
  OAI2BB2XL U1313 ( .B0(n1461), .B1(n1708), .A0N(\gbuff[15][28] ), .A1N(n1709), 
        .Y(n2310) );
  OAI2BB2XL U1314 ( .B0(n1459), .B1(n1708), .A0N(\gbuff[15][29] ), .A1N(n1709), 
        .Y(n2309) );
  OAI2BB2XL U1315 ( .B0(n1457), .B1(n1708), .A0N(\gbuff[15][30] ), .A1N(n1709), 
        .Y(n2308) );
  OAI2BB2XL U1316 ( .B0(n1455), .B1(n1708), .A0N(\gbuff[15][31] ), .A1N(n1707), 
        .Y(n2307) );
  OAI2BB2XL U1317 ( .B0(n1517), .B1(n1704), .A0N(\gbuff[16][0] ), .A1N(n1706), 
        .Y(n2306) );
  OAI2BB2XL U1318 ( .B0(n1515), .B1(n1704), .A0N(\gbuff[16][1] ), .A1N(n1705), 
        .Y(n2305) );
  OAI2BB2XL U1319 ( .B0(n1513), .B1(n1704), .A0N(\gbuff[16][2] ), .A1N(n1704), 
        .Y(n2304) );
  OAI2BB2XL U1320 ( .B0(n1511), .B1(n1704), .A0N(\gbuff[16][3] ), .A1N(n1706), 
        .Y(n2303) );
  OAI2BB2XL U1321 ( .B0(n1509), .B1(n1704), .A0N(\gbuff[16][4] ), .A1N(n1706), 
        .Y(n2302) );
  OAI2BB2XL U1322 ( .B0(n1507), .B1(n1704), .A0N(\gbuff[16][5] ), .A1N(n1706), 
        .Y(n2301) );
  OAI2BB2XL U1323 ( .B0(n1505), .B1(n1704), .A0N(\gbuff[16][6] ), .A1N(n1706), 
        .Y(n2300) );
  OAI2BB2XL U1324 ( .B0(n1503), .B1(n1704), .A0N(\gbuff[16][7] ), .A1N(n1706), 
        .Y(n2299) );
  OAI2BB2XL U1325 ( .B0(n1501), .B1(n1704), .A0N(\gbuff[16][8] ), .A1N(n1706), 
        .Y(n2298) );
  OAI2BB2XL U1326 ( .B0(n1499), .B1(n1704), .A0N(\gbuff[16][9] ), .A1N(n1706), 
        .Y(n2297) );
  OAI2BB2XL U1327 ( .B0(n1497), .B1(n1704), .A0N(\gbuff[16][10] ), .A1N(n1706), 
        .Y(n2296) );
  OAI2BB2XL U1328 ( .B0(n1495), .B1(n1704), .A0N(\gbuff[16][11] ), .A1N(n1706), 
        .Y(n2295) );
  OAI2BB2XL U1329 ( .B0(n1493), .B1(n1704), .A0N(\gbuff[16][12] ), .A1N(n1706), 
        .Y(n2294) );
  OAI2BB2XL U1330 ( .B0(n1491), .B1(n1704), .A0N(\gbuff[16][13] ), .A1N(n1706), 
        .Y(n2293) );
  OAI2BB2XL U1331 ( .B0(n1489), .B1(n1705), .A0N(\gbuff[16][14] ), .A1N(n1706), 
        .Y(n2292) );
  OAI2BB2XL U1332 ( .B0(n1487), .B1(n1704), .A0N(\gbuff[16][15] ), .A1N(n1705), 
        .Y(n2291) );
  OAI2BB2XL U1333 ( .B0(n1485), .B1(n1705), .A0N(\gbuff[16][16] ), .A1N(n1706), 
        .Y(n2290) );
  OAI2BB2XL U1334 ( .B0(n1483), .B1(n1704), .A0N(\gbuff[16][17] ), .A1N(n1705), 
        .Y(n2289) );
  OAI2BB2XL U1335 ( .B0(n1481), .B1(n1705), .A0N(\gbuff[16][18] ), .A1N(n1705), 
        .Y(n2288) );
  OAI2BB2XL U1336 ( .B0(n1479), .B1(n1704), .A0N(\gbuff[16][19] ), .A1N(n1705), 
        .Y(n2287) );
  OAI2BB2XL U1337 ( .B0(n1477), .B1(n1705), .A0N(\gbuff[16][20] ), .A1N(n1705), 
        .Y(n2286) );
  OAI2BB2XL U1338 ( .B0(n1475), .B1(n1704), .A0N(\gbuff[16][21] ), .A1N(n1705), 
        .Y(n2285) );
  OAI2BB2XL U1339 ( .B0(n1473), .B1(n1705), .A0N(\gbuff[16][22] ), .A1N(n1706), 
        .Y(n2284) );
  OAI2BB2XL U1340 ( .B0(n1471), .B1(n1705), .A0N(\gbuff[16][23] ), .A1N(n1705), 
        .Y(n2283) );
  OAI2BB2XL U1341 ( .B0(n1469), .B1(n1704), .A0N(\gbuff[16][24] ), .A1N(n1706), 
        .Y(n2282) );
  OAI2BB2XL U1342 ( .B0(n1467), .B1(n1705), .A0N(\gbuff[16][25] ), .A1N(n1706), 
        .Y(n2281) );
  OAI2BB2XL U1343 ( .B0(n1465), .B1(n1705), .A0N(\gbuff[16][26] ), .A1N(n1706), 
        .Y(n2280) );
  OAI2BB2XL U1344 ( .B0(n1463), .B1(n1705), .A0N(\gbuff[16][27] ), .A1N(n1706), 
        .Y(n2279) );
  OAI2BB2XL U1345 ( .B0(n1461), .B1(n1705), .A0N(\gbuff[16][28] ), .A1N(n1706), 
        .Y(n2278) );
  OAI2BB2XL U1346 ( .B0(n1459), .B1(n1705), .A0N(\gbuff[16][29] ), .A1N(n1706), 
        .Y(n2277) );
  OAI2BB2XL U1347 ( .B0(n1457), .B1(n1705), .A0N(\gbuff[16][30] ), .A1N(n1706), 
        .Y(n2276) );
  OAI2BB2XL U1348 ( .B0(n1455), .B1(n1705), .A0N(\gbuff[16][31] ), .A1N(n1704), 
        .Y(n2275) );
  OAI2BB2XL U1349 ( .B0(n1517), .B1(n1701), .A0N(\gbuff[17][0] ), .A1N(n1703), 
        .Y(n2274) );
  OAI2BB2XL U1350 ( .B0(n1515), .B1(n1701), .A0N(\gbuff[17][1] ), .A1N(n1702), 
        .Y(n2273) );
  OAI2BB2XL U1351 ( .B0(n1513), .B1(n1701), .A0N(\gbuff[17][2] ), .A1N(n1701), 
        .Y(n2272) );
  OAI2BB2XL U1352 ( .B0(n1511), .B1(n1701), .A0N(\gbuff[17][3] ), .A1N(n1703), 
        .Y(n2271) );
  OAI2BB2XL U1353 ( .B0(n1509), .B1(n1701), .A0N(\gbuff[17][4] ), .A1N(n1703), 
        .Y(n2270) );
  OAI2BB2XL U1354 ( .B0(n1507), .B1(n1701), .A0N(\gbuff[17][5] ), .A1N(n1703), 
        .Y(n2269) );
  OAI2BB2XL U1355 ( .B0(n1505), .B1(n1701), .A0N(\gbuff[17][6] ), .A1N(n1703), 
        .Y(n2268) );
  OAI2BB2XL U1356 ( .B0(n1503), .B1(n1701), .A0N(\gbuff[17][7] ), .A1N(n1703), 
        .Y(n2267) );
  OAI2BB2XL U1357 ( .B0(n1501), .B1(n1701), .A0N(\gbuff[17][8] ), .A1N(n1703), 
        .Y(n2266) );
  OAI2BB2XL U1358 ( .B0(n1499), .B1(n1701), .A0N(\gbuff[17][9] ), .A1N(n1703), 
        .Y(n2265) );
  OAI2BB2XL U1359 ( .B0(n1497), .B1(n1701), .A0N(\gbuff[17][10] ), .A1N(n1703), 
        .Y(n2264) );
  OAI2BB2XL U1360 ( .B0(n1495), .B1(n1701), .A0N(\gbuff[17][11] ), .A1N(n1703), 
        .Y(n2263) );
  OAI2BB2XL U1361 ( .B0(n1493), .B1(n1701), .A0N(\gbuff[17][12] ), .A1N(n1703), 
        .Y(n2262) );
  OAI2BB2XL U1362 ( .B0(n1491), .B1(n1701), .A0N(\gbuff[17][13] ), .A1N(n1703), 
        .Y(n2261) );
  OAI2BB2XL U1363 ( .B0(n1489), .B1(n1702), .A0N(\gbuff[17][14] ), .A1N(n1703), 
        .Y(n2260) );
  OAI2BB2XL U1364 ( .B0(n1487), .B1(n1701), .A0N(\gbuff[17][15] ), .A1N(n1702), 
        .Y(n2259) );
  OAI2BB2XL U1365 ( .B0(n1485), .B1(n1702), .A0N(\gbuff[17][16] ), .A1N(n1703), 
        .Y(n2258) );
  OAI2BB2XL U1366 ( .B0(n1483), .B1(n1701), .A0N(\gbuff[17][17] ), .A1N(n1702), 
        .Y(n2257) );
  OAI2BB2XL U1367 ( .B0(n1481), .B1(n1702), .A0N(\gbuff[17][18] ), .A1N(n1702), 
        .Y(n2256) );
  OAI2BB2XL U1368 ( .B0(n1479), .B1(n1701), .A0N(\gbuff[17][19] ), .A1N(n1702), 
        .Y(n2255) );
  OAI2BB2XL U1369 ( .B0(n1477), .B1(n1702), .A0N(\gbuff[17][20] ), .A1N(n1702), 
        .Y(n2254) );
  OAI2BB2XL U1370 ( .B0(n1475), .B1(n1701), .A0N(\gbuff[17][21] ), .A1N(n1702), 
        .Y(n2253) );
  OAI2BB2XL U1371 ( .B0(n1473), .B1(n1702), .A0N(\gbuff[17][22] ), .A1N(n1703), 
        .Y(n2252) );
  OAI2BB2XL U1372 ( .B0(n1471), .B1(n1702), .A0N(\gbuff[17][23] ), .A1N(n1702), 
        .Y(n2251) );
  OAI2BB2XL U1373 ( .B0(n1469), .B1(n1701), .A0N(\gbuff[17][24] ), .A1N(n1703), 
        .Y(n2250) );
  OAI2BB2XL U1374 ( .B0(n1467), .B1(n1702), .A0N(\gbuff[17][25] ), .A1N(n1703), 
        .Y(n2249) );
  OAI2BB2XL U1375 ( .B0(n1465), .B1(n1702), .A0N(\gbuff[17][26] ), .A1N(n1703), 
        .Y(n2248) );
  OAI2BB2XL U1376 ( .B0(n1463), .B1(n1702), .A0N(\gbuff[17][27] ), .A1N(n1703), 
        .Y(n2247) );
  OAI2BB2XL U1377 ( .B0(n1461), .B1(n1702), .A0N(\gbuff[17][28] ), .A1N(n1703), 
        .Y(n2246) );
  OAI2BB2XL U1378 ( .B0(n1459), .B1(n1702), .A0N(\gbuff[17][29] ), .A1N(n1703), 
        .Y(n2245) );
  OAI2BB2XL U1379 ( .B0(n1457), .B1(n1702), .A0N(\gbuff[17][30] ), .A1N(n1703), 
        .Y(n2244) );
  OAI2BB2XL U1380 ( .B0(n1455), .B1(n1702), .A0N(\gbuff[17][31] ), .A1N(n1701), 
        .Y(n2243) );
  OAI2BB2XL U1381 ( .B0(n1517), .B1(n1698), .A0N(\gbuff[18][0] ), .A1N(n1700), 
        .Y(n2242) );
  OAI2BB2XL U1382 ( .B0(n1515), .B1(n1698), .A0N(\gbuff[18][1] ), .A1N(n1699), 
        .Y(n2241) );
  OAI2BB2XL U1383 ( .B0(n1513), .B1(n1698), .A0N(\gbuff[18][2] ), .A1N(n1698), 
        .Y(n2240) );
  OAI2BB2XL U1384 ( .B0(n1511), .B1(n1698), .A0N(\gbuff[18][3] ), .A1N(n1700), 
        .Y(n2239) );
  OAI2BB2XL U1385 ( .B0(n1509), .B1(n1698), .A0N(\gbuff[18][4] ), .A1N(n1700), 
        .Y(n2238) );
  OAI2BB2XL U1386 ( .B0(n1507), .B1(n1698), .A0N(\gbuff[18][5] ), .A1N(n1700), 
        .Y(n2237) );
  OAI2BB2XL U1387 ( .B0(n1505), .B1(n1698), .A0N(\gbuff[18][6] ), .A1N(n1700), 
        .Y(n2236) );
  OAI2BB2XL U1388 ( .B0(n1503), .B1(n1698), .A0N(\gbuff[18][7] ), .A1N(n1700), 
        .Y(n2235) );
  OAI2BB2XL U1389 ( .B0(n1501), .B1(n1698), .A0N(\gbuff[18][8] ), .A1N(n1700), 
        .Y(n2234) );
  OAI2BB2XL U1390 ( .B0(n1499), .B1(n1698), .A0N(\gbuff[18][9] ), .A1N(n1700), 
        .Y(n2233) );
  OAI2BB2XL U1391 ( .B0(n1497), .B1(n1698), .A0N(\gbuff[18][10] ), .A1N(n1700), 
        .Y(n2232) );
  OAI2BB2XL U1392 ( .B0(n1495), .B1(n1698), .A0N(\gbuff[18][11] ), .A1N(n1700), 
        .Y(n2231) );
  OAI2BB2XL U1393 ( .B0(n1493), .B1(n1698), .A0N(\gbuff[18][12] ), .A1N(n1700), 
        .Y(n2230) );
  OAI2BB2XL U1394 ( .B0(n1491), .B1(n1698), .A0N(\gbuff[18][13] ), .A1N(n1700), 
        .Y(n2229) );
  OAI2BB2XL U1395 ( .B0(n1489), .B1(n1699), .A0N(\gbuff[18][14] ), .A1N(n1700), 
        .Y(n2228) );
  OAI2BB2XL U1396 ( .B0(n1487), .B1(n1698), .A0N(\gbuff[18][15] ), .A1N(n1699), 
        .Y(n2227) );
  OAI2BB2XL U1397 ( .B0(n1485), .B1(n1699), .A0N(\gbuff[18][16] ), .A1N(n1700), 
        .Y(n2226) );
  OAI2BB2XL U1398 ( .B0(n1483), .B1(n1698), .A0N(\gbuff[18][17] ), .A1N(n1699), 
        .Y(n2225) );
  OAI2BB2XL U1399 ( .B0(n1481), .B1(n1699), .A0N(\gbuff[18][18] ), .A1N(n1699), 
        .Y(n2224) );
  OAI2BB2XL U1400 ( .B0(n1479), .B1(n1698), .A0N(\gbuff[18][19] ), .A1N(n1699), 
        .Y(n2223) );
  OAI2BB2XL U1401 ( .B0(n1477), .B1(n1699), .A0N(\gbuff[18][20] ), .A1N(n1699), 
        .Y(n2222) );
  OAI2BB2XL U1402 ( .B0(n1475), .B1(n1698), .A0N(\gbuff[18][21] ), .A1N(n1699), 
        .Y(n2221) );
  OAI2BB2XL U1403 ( .B0(n1473), .B1(n1699), .A0N(\gbuff[18][22] ), .A1N(n1700), 
        .Y(n2220) );
  OAI2BB2XL U1404 ( .B0(n1471), .B1(n1699), .A0N(\gbuff[18][23] ), .A1N(n1699), 
        .Y(n2219) );
  OAI2BB2XL U1405 ( .B0(n1469), .B1(n1698), .A0N(\gbuff[18][24] ), .A1N(n1700), 
        .Y(n2218) );
  OAI2BB2XL U1406 ( .B0(n1467), .B1(n1699), .A0N(\gbuff[18][25] ), .A1N(n1700), 
        .Y(n2217) );
  OAI2BB2XL U1407 ( .B0(n1465), .B1(n1699), .A0N(\gbuff[18][26] ), .A1N(n1700), 
        .Y(n2216) );
  OAI2BB2XL U1408 ( .B0(n1463), .B1(n1699), .A0N(\gbuff[18][27] ), .A1N(n1700), 
        .Y(n2215) );
  OAI2BB2XL U1409 ( .B0(n1461), .B1(n1699), .A0N(\gbuff[18][28] ), .A1N(n1700), 
        .Y(n2214) );
  OAI2BB2XL U1410 ( .B0(n1459), .B1(n1699), .A0N(\gbuff[18][29] ), .A1N(n1700), 
        .Y(n2213) );
  OAI2BB2XL U1411 ( .B0(n1457), .B1(n1699), .A0N(\gbuff[18][30] ), .A1N(n1700), 
        .Y(n2212) );
  OAI2BB2XL U1412 ( .B0(n1455), .B1(n1699), .A0N(\gbuff[18][31] ), .A1N(n1698), 
        .Y(n2211) );
  OAI2BB2XL U1413 ( .B0(n1517), .B1(n1695), .A0N(\gbuff[19][0] ), .A1N(n1697), 
        .Y(n2210) );
  OAI2BB2XL U1414 ( .B0(n1515), .B1(n1695), .A0N(\gbuff[19][1] ), .A1N(n1696), 
        .Y(n2209) );
  OAI2BB2XL U1415 ( .B0(n1513), .B1(n1695), .A0N(\gbuff[19][2] ), .A1N(n1695), 
        .Y(n2208) );
  OAI2BB2XL U1416 ( .B0(n1511), .B1(n1695), .A0N(\gbuff[19][3] ), .A1N(n1697), 
        .Y(n2207) );
  OAI2BB2XL U1417 ( .B0(n1509), .B1(n1695), .A0N(\gbuff[19][4] ), .A1N(n1697), 
        .Y(n2206) );
  OAI2BB2XL U1418 ( .B0(n1507), .B1(n1695), .A0N(\gbuff[19][5] ), .A1N(n1697), 
        .Y(n2205) );
  OAI2BB2XL U1419 ( .B0(n1505), .B1(n1695), .A0N(\gbuff[19][6] ), .A1N(n1697), 
        .Y(n2204) );
  OAI2BB2XL U1420 ( .B0(n1503), .B1(n1695), .A0N(\gbuff[19][7] ), .A1N(n1697), 
        .Y(n2203) );
  OAI2BB2XL U1421 ( .B0(n1501), .B1(n1695), .A0N(\gbuff[19][8] ), .A1N(n1697), 
        .Y(n2202) );
  OAI2BB2XL U1422 ( .B0(n1499), .B1(n1695), .A0N(\gbuff[19][9] ), .A1N(n1697), 
        .Y(n2201) );
  OAI2BB2XL U1423 ( .B0(n1497), .B1(n1695), .A0N(\gbuff[19][10] ), .A1N(n1697), 
        .Y(n2200) );
  OAI2BB2XL U1424 ( .B0(n1495), .B1(n1695), .A0N(\gbuff[19][11] ), .A1N(n1697), 
        .Y(n2199) );
  OAI2BB2XL U1425 ( .B0(n1493), .B1(n1695), .A0N(\gbuff[19][12] ), .A1N(n1697), 
        .Y(n2198) );
  OAI2BB2XL U1426 ( .B0(n1491), .B1(n1695), .A0N(\gbuff[19][13] ), .A1N(n1697), 
        .Y(n2197) );
  OAI2BB2XL U1427 ( .B0(n1489), .B1(n1696), .A0N(\gbuff[19][14] ), .A1N(n1697), 
        .Y(n2196) );
  OAI2BB2XL U1428 ( .B0(n1487), .B1(n1695), .A0N(\gbuff[19][15] ), .A1N(n1696), 
        .Y(n2195) );
  OAI2BB2XL U1429 ( .B0(n1485), .B1(n1696), .A0N(\gbuff[19][16] ), .A1N(n1697), 
        .Y(n2194) );
  OAI2BB2XL U1430 ( .B0(n1483), .B1(n1695), .A0N(\gbuff[19][17] ), .A1N(n1696), 
        .Y(n2193) );
  OAI2BB2XL U1431 ( .B0(n1481), .B1(n1696), .A0N(\gbuff[19][18] ), .A1N(n1696), 
        .Y(n2192) );
  OAI2BB2XL U1432 ( .B0(n1479), .B1(n1695), .A0N(\gbuff[19][19] ), .A1N(n1696), 
        .Y(n2191) );
  OAI2BB2XL U1433 ( .B0(n1477), .B1(n1696), .A0N(\gbuff[19][20] ), .A1N(n1696), 
        .Y(n2190) );
  OAI2BB2XL U1434 ( .B0(n1475), .B1(n1695), .A0N(\gbuff[19][21] ), .A1N(n1696), 
        .Y(n2189) );
  OAI2BB2XL U1435 ( .B0(n1473), .B1(n1696), .A0N(\gbuff[19][22] ), .A1N(n1697), 
        .Y(n2188) );
  OAI2BB2XL U1436 ( .B0(n1471), .B1(n1696), .A0N(\gbuff[19][23] ), .A1N(n1696), 
        .Y(n2187) );
  OAI2BB2XL U1437 ( .B0(n1469), .B1(n1695), .A0N(\gbuff[19][24] ), .A1N(n1697), 
        .Y(n2186) );
  OAI2BB2XL U1438 ( .B0(n1467), .B1(n1696), .A0N(\gbuff[19][25] ), .A1N(n1697), 
        .Y(n2185) );
  OAI2BB2XL U1439 ( .B0(n1465), .B1(n1696), .A0N(\gbuff[19][26] ), .A1N(n1697), 
        .Y(n2184) );
  OAI2BB2XL U1440 ( .B0(n1463), .B1(n1696), .A0N(\gbuff[19][27] ), .A1N(n1697), 
        .Y(n2183) );
  OAI2BB2XL U1441 ( .B0(n1461), .B1(n1696), .A0N(\gbuff[19][28] ), .A1N(n1697), 
        .Y(n2182) );
  OAI2BB2XL U1442 ( .B0(n1459), .B1(n1696), .A0N(\gbuff[19][29] ), .A1N(n1697), 
        .Y(n2181) );
  OAI2BB2XL U1443 ( .B0(n1457), .B1(n1696), .A0N(\gbuff[19][30] ), .A1N(n1697), 
        .Y(n2180) );
  OAI2BB2XL U1444 ( .B0(n1455), .B1(n1696), .A0N(\gbuff[19][31] ), .A1N(n1695), 
        .Y(n2179) );
  OAI2BB2XL U1445 ( .B0(n1516), .B1(n1692), .A0N(\gbuff[20][0] ), .A1N(n1693), 
        .Y(n2178) );
  OAI2BB2XL U1446 ( .B0(n1514), .B1(n1692), .A0N(\gbuff[20][1] ), .A1N(n1692), 
        .Y(n2177) );
  OAI2BB2XL U1447 ( .B0(n1512), .B1(n1692), .A0N(\gbuff[20][2] ), .A1N(n1694), 
        .Y(n2176) );
  OAI2BB2XL U1448 ( .B0(n1510), .B1(n1692), .A0N(\gbuff[20][3] ), .A1N(n1694), 
        .Y(n2175) );
  OAI2BB2XL U1449 ( .B0(n1508), .B1(n1692), .A0N(\gbuff[20][4] ), .A1N(n1692), 
        .Y(n2174) );
  OAI2BB2XL U1450 ( .B0(n1506), .B1(n1692), .A0N(\gbuff[20][5] ), .A1N(n1694), 
        .Y(n2173) );
  OAI2BB2XL U1451 ( .B0(n1504), .B1(n1692), .A0N(\gbuff[20][6] ), .A1N(n1694), 
        .Y(n2172) );
  OAI2BB2XL U1452 ( .B0(n1502), .B1(n1692), .A0N(\gbuff[20][7] ), .A1N(n1694), 
        .Y(n2171) );
  OAI2BB2XL U1453 ( .B0(n1500), .B1(n1692), .A0N(\gbuff[20][8] ), .A1N(n1694), 
        .Y(n2170) );
  OAI2BB2XL U1454 ( .B0(n1498), .B1(n1692), .A0N(\gbuff[20][9] ), .A1N(n1694), 
        .Y(n2169) );
  OAI2BB2XL U1455 ( .B0(n1496), .B1(n1692), .A0N(\gbuff[20][10] ), .A1N(n1694), 
        .Y(n2168) );
  OAI2BB2XL U1456 ( .B0(n1494), .B1(n1692), .A0N(\gbuff[20][11] ), .A1N(n1694), 
        .Y(n2167) );
  OAI2BB2XL U1457 ( .B0(n1492), .B1(n1692), .A0N(\gbuff[20][12] ), .A1N(n1694), 
        .Y(n2166) );
  OAI2BB2XL U1458 ( .B0(n1490), .B1(n1692), .A0N(\gbuff[20][13] ), .A1N(n1694), 
        .Y(n2165) );
  OAI2BB2XL U1459 ( .B0(n1488), .B1(n1692), .A0N(\gbuff[20][14] ), .A1N(n1694), 
        .Y(n2164) );
  OAI2BB2XL U1460 ( .B0(n1486), .B1(n1692), .A0N(\gbuff[20][15] ), .A1N(n1693), 
        .Y(n2163) );
  OAI2BB2XL U1461 ( .B0(n1484), .B1(n1692), .A0N(\gbuff[20][16] ), .A1N(n1694), 
        .Y(n2162) );
  OAI2BB2XL U1462 ( .B0(n1482), .B1(n1693), .A0N(\gbuff[20][17] ), .A1N(n1693), 
        .Y(n2161) );
  OAI2BB2XL U1463 ( .B0(n1480), .B1(n1692), .A0N(\gbuff[20][18] ), .A1N(n1693), 
        .Y(n2160) );
  OAI2BB2XL U1464 ( .B0(n1478), .B1(n1693), .A0N(\gbuff[20][19] ), .A1N(n1693), 
        .Y(n2159) );
  OAI2BB2XL U1465 ( .B0(n1476), .B1(n1692), .A0N(\gbuff[20][20] ), .A1N(n1693), 
        .Y(n2158) );
  OAI2BB2XL U1466 ( .B0(n1474), .B1(n1693), .A0N(\gbuff[20][21] ), .A1N(n1693), 
        .Y(n2157) );
  OAI2BB2XL U1467 ( .B0(n1472), .B1(n1693), .A0N(\gbuff[20][22] ), .A1N(n1694), 
        .Y(n2156) );
  OAI2BB2XL U1468 ( .B0(n1470), .B1(n1693), .A0N(\gbuff[20][23] ), .A1N(n1693), 
        .Y(n2155) );
  OAI2BB2XL U1469 ( .B0(n1468), .B1(n1694), .A0N(\gbuff[20][24] ), .A1N(n1694), 
        .Y(n2154) );
  OAI2BB2XL U1470 ( .B0(n1466), .B1(n1693), .A0N(\gbuff[20][25] ), .A1N(n1694), 
        .Y(n2153) );
  OAI2BB2XL U1471 ( .B0(n1464), .B1(n1693), .A0N(\gbuff[20][26] ), .A1N(n1694), 
        .Y(n2152) );
  OAI2BB2XL U1472 ( .B0(n1462), .B1(n1693), .A0N(\gbuff[20][27] ), .A1N(n1694), 
        .Y(n2151) );
  OAI2BB2XL U1473 ( .B0(n1460), .B1(n1693), .A0N(\gbuff[20][28] ), .A1N(n1694), 
        .Y(n2150) );
  OAI2BB2XL U1474 ( .B0(n1458), .B1(n1693), .A0N(\gbuff[20][29] ), .A1N(n1694), 
        .Y(n2149) );
  OAI2BB2XL U1475 ( .B0(n1456), .B1(n1693), .A0N(\gbuff[20][30] ), .A1N(n2831), 
        .Y(n2148) );
  OAI2BB2XL U1476 ( .B0(n1454), .B1(n1693), .A0N(\gbuff[20][31] ), .A1N(n2831), 
        .Y(n2147) );
  OAI2BB2XL U1477 ( .B0(n1516), .B1(n1689), .A0N(\gbuff[21][0] ), .A1N(n1691), 
        .Y(n2146) );
  OAI2BB2XL U1478 ( .B0(n1514), .B1(n1689), .A0N(\gbuff[21][1] ), .A1N(n2830), 
        .Y(n2145) );
  OAI2BB2XL U1479 ( .B0(n1512), .B1(n1689), .A0N(\gbuff[21][2] ), .A1N(n1689), 
        .Y(n2144) );
  OAI2BB2XL U1480 ( .B0(n1510), .B1(n1689), .A0N(\gbuff[21][3] ), .A1N(n1691), 
        .Y(n2143) );
  OAI2BB2XL U1481 ( .B0(n1508), .B1(n1689), .A0N(\gbuff[21][4] ), .A1N(n1691), 
        .Y(n2142) );
  OAI2BB2XL U1482 ( .B0(n1506), .B1(n1689), .A0N(\gbuff[21][5] ), .A1N(n1691), 
        .Y(n2141) );
  OAI2BB2XL U1483 ( .B0(n1504), .B1(n1689), .A0N(\gbuff[21][6] ), .A1N(n1691), 
        .Y(n2140) );
  OAI2BB2XL U1484 ( .B0(n1502), .B1(n1689), .A0N(\gbuff[21][7] ), .A1N(n1691), 
        .Y(n2139) );
  OAI2BB2XL U1485 ( .B0(n1500), .B1(n1689), .A0N(\gbuff[21][8] ), .A1N(n1691), 
        .Y(n2138) );
  OAI2BB2XL U1486 ( .B0(n1498), .B1(n1689), .A0N(\gbuff[21][9] ), .A1N(n1691), 
        .Y(n2137) );
  OAI2BB2XL U1487 ( .B0(n1496), .B1(n1689), .A0N(\gbuff[21][10] ), .A1N(n1691), 
        .Y(n2136) );
  OAI2BB2XL U1488 ( .B0(n1494), .B1(n1689), .A0N(\gbuff[21][11] ), .A1N(n1691), 
        .Y(n2135) );
  OAI2BB2XL U1489 ( .B0(n1492), .B1(n1689), .A0N(\gbuff[21][12] ), .A1N(n1691), 
        .Y(n2134) );
  OAI2BB2XL U1490 ( .B0(n1490), .B1(n1689), .A0N(\gbuff[21][13] ), .A1N(n1691), 
        .Y(n2133) );
  OAI2BB2XL U1491 ( .B0(n1488), .B1(n1690), .A0N(\gbuff[21][14] ), .A1N(n1691), 
        .Y(n2132) );
  OAI2BB2XL U1492 ( .B0(n1486), .B1(n1689), .A0N(\gbuff[21][15] ), .A1N(n1690), 
        .Y(n2131) );
  OAI2BB2XL U1493 ( .B0(n1484), .B1(n1690), .A0N(\gbuff[21][16] ), .A1N(n1691), 
        .Y(n2130) );
  OAI2BB2XL U1494 ( .B0(n1482), .B1(n1689), .A0N(\gbuff[21][17] ), .A1N(n1690), 
        .Y(n2129) );
  OAI2BB2XL U1495 ( .B0(n1480), .B1(n1690), .A0N(\gbuff[21][18] ), .A1N(n1690), 
        .Y(n2128) );
  OAI2BB2XL U1496 ( .B0(n1478), .B1(n1689), .A0N(\gbuff[21][19] ), .A1N(n1690), 
        .Y(n2127) );
  OAI2BB2XL U1497 ( .B0(n1476), .B1(n1690), .A0N(\gbuff[21][20] ), .A1N(n1690), 
        .Y(n2126) );
  OAI2BB2XL U1498 ( .B0(n1474), .B1(n1689), .A0N(\gbuff[21][21] ), .A1N(n1690), 
        .Y(n2125) );
  OAI2BB2XL U1499 ( .B0(n1472), .B1(n1690), .A0N(\gbuff[21][22] ), .A1N(n1691), 
        .Y(n2124) );
  OAI2BB2XL U1500 ( .B0(n1470), .B1(n1690), .A0N(\gbuff[21][23] ), .A1N(n1690), 
        .Y(n2123) );
  OAI2BB2XL U1501 ( .B0(n1468), .B1(n2830), .A0N(\gbuff[21][24] ), .A1N(n1691), 
        .Y(n2122) );
  OAI2BB2XL U1502 ( .B0(n1466), .B1(n1690), .A0N(\gbuff[21][25] ), .A1N(n1691), 
        .Y(n2121) );
  OAI2BB2XL U1503 ( .B0(n1464), .B1(n1690), .A0N(\gbuff[21][26] ), .A1N(n1691), 
        .Y(n2120) );
  OAI2BB2XL U1504 ( .B0(n1462), .B1(n1690), .A0N(\gbuff[21][27] ), .A1N(n1691), 
        .Y(n2119) );
  OAI2BB2XL U1505 ( .B0(n1460), .B1(n1690), .A0N(\gbuff[21][28] ), .A1N(n1691), 
        .Y(n2118) );
  OAI2BB2XL U1506 ( .B0(n1458), .B1(n1690), .A0N(\gbuff[21][29] ), .A1N(n1691), 
        .Y(n2117) );
  OAI2BB2XL U1507 ( .B0(n1456), .B1(n1690), .A0N(\gbuff[21][30] ), .A1N(n1691), 
        .Y(n2116) );
  OAI2BB2XL U1508 ( .B0(n1454), .B1(n1690), .A0N(\gbuff[21][31] ), .A1N(n1689), 
        .Y(n2115) );
  OAI2BB2XL U1509 ( .B0(n1516), .B1(n1686), .A0N(\gbuff[22][0] ), .A1N(n1688), 
        .Y(n2114) );
  OAI2BB2XL U1510 ( .B0(n1514), .B1(n1686), .A0N(\gbuff[22][1] ), .A1N(n2829), 
        .Y(n2113) );
  OAI2BB2XL U1511 ( .B0(n1512), .B1(n1686), .A0N(\gbuff[22][2] ), .A1N(n1686), 
        .Y(n2112) );
  OAI2BB2XL U1512 ( .B0(n1510), .B1(n1686), .A0N(\gbuff[22][3] ), .A1N(n1688), 
        .Y(n2111) );
  OAI2BB2XL U1513 ( .B0(n1508), .B1(n1686), .A0N(\gbuff[22][4] ), .A1N(n1688), 
        .Y(n2110) );
  OAI2BB2XL U1514 ( .B0(n1506), .B1(n1686), .A0N(\gbuff[22][5] ), .A1N(n1688), 
        .Y(n2109) );
  OAI2BB2XL U1515 ( .B0(n1504), .B1(n1686), .A0N(\gbuff[22][6] ), .A1N(n1688), 
        .Y(n2108) );
  OAI2BB2XL U1516 ( .B0(n1502), .B1(n1686), .A0N(\gbuff[22][7] ), .A1N(n1688), 
        .Y(n2107) );
  OAI2BB2XL U1517 ( .B0(n1500), .B1(n1686), .A0N(\gbuff[22][8] ), .A1N(n1688), 
        .Y(n2106) );
  OAI2BB2XL U1518 ( .B0(n1498), .B1(n1686), .A0N(\gbuff[22][9] ), .A1N(n1688), 
        .Y(n2105) );
  OAI2BB2XL U1519 ( .B0(n1496), .B1(n1686), .A0N(\gbuff[22][10] ), .A1N(n1688), 
        .Y(n2104) );
  OAI2BB2XL U1520 ( .B0(n1494), .B1(n1686), .A0N(\gbuff[22][11] ), .A1N(n1688), 
        .Y(n2103) );
  OAI2BB2XL U1521 ( .B0(n1492), .B1(n1686), .A0N(\gbuff[22][12] ), .A1N(n1688), 
        .Y(n2102) );
  OAI2BB2XL U1522 ( .B0(n1490), .B1(n1686), .A0N(\gbuff[22][13] ), .A1N(n1688), 
        .Y(n2101) );
  OAI2BB2XL U1523 ( .B0(n1488), .B1(n1687), .A0N(\gbuff[22][14] ), .A1N(n1688), 
        .Y(n2100) );
  OAI2BB2XL U1524 ( .B0(n1486), .B1(n1686), .A0N(\gbuff[22][15] ), .A1N(n1687), 
        .Y(n2099) );
  OAI2BB2XL U1525 ( .B0(n1484), .B1(n1687), .A0N(\gbuff[22][16] ), .A1N(n1688), 
        .Y(n2098) );
  OAI2BB2XL U1526 ( .B0(n1482), .B1(n1686), .A0N(\gbuff[22][17] ), .A1N(n1687), 
        .Y(n2097) );
  OAI2BB2XL U1527 ( .B0(n1480), .B1(n1687), .A0N(\gbuff[22][18] ), .A1N(n1687), 
        .Y(n2096) );
  OAI2BB2XL U1528 ( .B0(n1478), .B1(n1686), .A0N(\gbuff[22][19] ), .A1N(n1687), 
        .Y(n2095) );
  OAI2BB2XL U1529 ( .B0(n1476), .B1(n1687), .A0N(\gbuff[22][20] ), .A1N(n1687), 
        .Y(n2094) );
  OAI2BB2XL U1530 ( .B0(n1474), .B1(n1686), .A0N(\gbuff[22][21] ), .A1N(n1687), 
        .Y(n2093) );
  OAI2BB2XL U1531 ( .B0(n1472), .B1(n1687), .A0N(\gbuff[22][22] ), .A1N(n1688), 
        .Y(n2092) );
  OAI2BB2XL U1532 ( .B0(n1470), .B1(n1687), .A0N(\gbuff[22][23] ), .A1N(n1687), 
        .Y(n2091) );
  OAI2BB2XL U1533 ( .B0(n1468), .B1(n2829), .A0N(\gbuff[22][24] ), .A1N(n1688), 
        .Y(n2090) );
  OAI2BB2XL U1534 ( .B0(n1466), .B1(n1687), .A0N(\gbuff[22][25] ), .A1N(n1688), 
        .Y(n2089) );
  OAI2BB2XL U1535 ( .B0(n1464), .B1(n1687), .A0N(\gbuff[22][26] ), .A1N(n1688), 
        .Y(n2088) );
  OAI2BB2XL U1536 ( .B0(n1462), .B1(n1687), .A0N(\gbuff[22][27] ), .A1N(n1688), 
        .Y(n2087) );
  OAI2BB2XL U1537 ( .B0(n1460), .B1(n1687), .A0N(\gbuff[22][28] ), .A1N(n1688), 
        .Y(n2086) );
  OAI2BB2XL U1538 ( .B0(n1458), .B1(n1687), .A0N(\gbuff[22][29] ), .A1N(n1688), 
        .Y(n2085) );
  OAI2BB2XL U1539 ( .B0(n1456), .B1(n1687), .A0N(\gbuff[22][30] ), .A1N(n1688), 
        .Y(n2084) );
  OAI2BB2XL U1540 ( .B0(n1454), .B1(n1687), .A0N(\gbuff[22][31] ), .A1N(n1686), 
        .Y(n2083) );
  OAI2BB2XL U1541 ( .B0(n1516), .B1(n1683), .A0N(\gbuff[23][0] ), .A1N(n1685), 
        .Y(n2082) );
  OAI2BB2XL U1542 ( .B0(n1514), .B1(n1683), .A0N(\gbuff[23][1] ), .A1N(n2828), 
        .Y(n2081) );
  OAI2BB2XL U1543 ( .B0(n1512), .B1(n1683), .A0N(\gbuff[23][2] ), .A1N(n1683), 
        .Y(n2080) );
  OAI2BB2XL U1544 ( .B0(n1510), .B1(n1683), .A0N(\gbuff[23][3] ), .A1N(n1685), 
        .Y(n2079) );
  OAI2BB2XL U1545 ( .B0(n1508), .B1(n1683), .A0N(\gbuff[23][4] ), .A1N(n1685), 
        .Y(n2078) );
  OAI2BB2XL U1546 ( .B0(n1506), .B1(n1683), .A0N(\gbuff[23][5] ), .A1N(n1685), 
        .Y(n2077) );
  OAI2BB2XL U1547 ( .B0(n1504), .B1(n1683), .A0N(\gbuff[23][6] ), .A1N(n1685), 
        .Y(n2076) );
  OAI2BB2XL U1548 ( .B0(n1502), .B1(n1683), .A0N(\gbuff[23][7] ), .A1N(n1685), 
        .Y(n2075) );
  OAI2BB2XL U1549 ( .B0(n1500), .B1(n1683), .A0N(\gbuff[23][8] ), .A1N(n1685), 
        .Y(n2074) );
  OAI2BB2XL U1550 ( .B0(n1498), .B1(n1683), .A0N(\gbuff[23][9] ), .A1N(n1685), 
        .Y(n2073) );
  OAI2BB2XL U1551 ( .B0(n1496), .B1(n1683), .A0N(\gbuff[23][10] ), .A1N(n1685), 
        .Y(n2072) );
  OAI2BB2XL U1552 ( .B0(n1494), .B1(n1683), .A0N(\gbuff[23][11] ), .A1N(n1685), 
        .Y(n2071) );
  OAI2BB2XL U1553 ( .B0(n1492), .B1(n1683), .A0N(\gbuff[23][12] ), .A1N(n1685), 
        .Y(n2070) );
  OAI2BB2XL U1554 ( .B0(n1490), .B1(n1683), .A0N(\gbuff[23][13] ), .A1N(n1685), 
        .Y(n2069) );
  OAI2BB2XL U1555 ( .B0(n1488), .B1(n1684), .A0N(\gbuff[23][14] ), .A1N(n1685), 
        .Y(n2068) );
  OAI2BB2XL U1556 ( .B0(n1486), .B1(n1683), .A0N(\gbuff[23][15] ), .A1N(n1684), 
        .Y(n2067) );
  OAI2BB2XL U1557 ( .B0(n1484), .B1(n1684), .A0N(\gbuff[23][16] ), .A1N(n1685), 
        .Y(n2066) );
  OAI2BB2XL U1558 ( .B0(n1482), .B1(n1683), .A0N(\gbuff[23][17] ), .A1N(n1684), 
        .Y(n2065) );
  OAI2BB2XL U1559 ( .B0(n1480), .B1(n1684), .A0N(\gbuff[23][18] ), .A1N(n1684), 
        .Y(n2064) );
  OAI2BB2XL U1560 ( .B0(n1478), .B1(n1683), .A0N(\gbuff[23][19] ), .A1N(n1684), 
        .Y(n2063) );
  OAI2BB2XL U1561 ( .B0(n1476), .B1(n1684), .A0N(\gbuff[23][20] ), .A1N(n1684), 
        .Y(n2062) );
  OAI2BB2XL U1562 ( .B0(n1474), .B1(n1683), .A0N(\gbuff[23][21] ), .A1N(n1684), 
        .Y(n2061) );
  OAI2BB2XL U1563 ( .B0(n1472), .B1(n1684), .A0N(\gbuff[23][22] ), .A1N(n1685), 
        .Y(n2060) );
  OAI2BB2XL U1564 ( .B0(n1470), .B1(n1684), .A0N(\gbuff[23][23] ), .A1N(n1684), 
        .Y(n2059) );
  OAI2BB2XL U1565 ( .B0(n1468), .B1(n2828), .A0N(\gbuff[23][24] ), .A1N(n1685), 
        .Y(n2058) );
  OAI2BB2XL U1566 ( .B0(n1466), .B1(n1684), .A0N(\gbuff[23][25] ), .A1N(n1685), 
        .Y(n2057) );
  OAI2BB2XL U1567 ( .B0(n1464), .B1(n1684), .A0N(\gbuff[23][26] ), .A1N(n1685), 
        .Y(n2056) );
  OAI2BB2XL U1568 ( .B0(n1462), .B1(n1684), .A0N(\gbuff[23][27] ), .A1N(n1685), 
        .Y(n2055) );
  OAI2BB2XL U1569 ( .B0(n1460), .B1(n1684), .A0N(\gbuff[23][28] ), .A1N(n1685), 
        .Y(n2054) );
  OAI2BB2XL U1570 ( .B0(n1458), .B1(n1684), .A0N(\gbuff[23][29] ), .A1N(n1685), 
        .Y(n2053) );
  OAI2BB2XL U1571 ( .B0(n1456), .B1(n1684), .A0N(\gbuff[23][30] ), .A1N(n1685), 
        .Y(n2052) );
  OAI2BB2XL U1572 ( .B0(n1454), .B1(n1684), .A0N(\gbuff[23][31] ), .A1N(n1683), 
        .Y(n2051) );
  OAI2BB2XL U1573 ( .B0(n1516), .B1(n1680), .A0N(\gbuff[24][0] ), .A1N(n1682), 
        .Y(n2050) );
  OAI2BB2XL U1574 ( .B0(n1514), .B1(n1680), .A0N(\gbuff[24][1] ), .A1N(n1681), 
        .Y(n2049) );
  OAI2BB2XL U1575 ( .B0(n1512), .B1(n1680), .A0N(\gbuff[24][2] ), .A1N(n1680), 
        .Y(n2048) );
  OAI2BB2XL U1576 ( .B0(n1510), .B1(n1680), .A0N(\gbuff[24][3] ), .A1N(n1682), 
        .Y(n2047) );
  OAI2BB2XL U1577 ( .B0(n1508), .B1(n1680), .A0N(\gbuff[24][4] ), .A1N(n1682), 
        .Y(n2046) );
  OAI2BB2XL U1578 ( .B0(n1506), .B1(n1680), .A0N(\gbuff[24][5] ), .A1N(n1682), 
        .Y(n2045) );
  OAI2BB2XL U1579 ( .B0(n1504), .B1(n1680), .A0N(\gbuff[24][6] ), .A1N(n1682), 
        .Y(n2044) );
  OAI2BB2XL U1580 ( .B0(n1502), .B1(n1680), .A0N(\gbuff[24][7] ), .A1N(n1682), 
        .Y(n2043) );
  OAI2BB2XL U1581 ( .B0(n1500), .B1(n1680), .A0N(\gbuff[24][8] ), .A1N(n1682), 
        .Y(n2042) );
  OAI2BB2XL U1582 ( .B0(n1498), .B1(n1680), .A0N(\gbuff[24][9] ), .A1N(n1682), 
        .Y(n2041) );
  OAI2BB2XL U1583 ( .B0(n1496), .B1(n1680), .A0N(\gbuff[24][10] ), .A1N(n1682), 
        .Y(n2040) );
  OAI2BB2XL U1584 ( .B0(n1494), .B1(n1680), .A0N(\gbuff[24][11] ), .A1N(n1682), 
        .Y(n2039) );
  OAI2BB2XL U1585 ( .B0(n1492), .B1(n1680), .A0N(\gbuff[24][12] ), .A1N(n1682), 
        .Y(n2038) );
  OAI2BB2XL U1586 ( .B0(n1490), .B1(n1680), .A0N(\gbuff[24][13] ), .A1N(n1682), 
        .Y(n2037) );
  OAI2BB2XL U1587 ( .B0(n1488), .B1(n1681), .A0N(\gbuff[24][14] ), .A1N(n1682), 
        .Y(n2036) );
  OAI2BB2XL U1588 ( .B0(n1486), .B1(n1680), .A0N(\gbuff[24][15] ), .A1N(n1681), 
        .Y(n2035) );
  OAI2BB2XL U1589 ( .B0(n1484), .B1(n1681), .A0N(\gbuff[24][16] ), .A1N(n1682), 
        .Y(n2034) );
  OAI2BB2XL U1590 ( .B0(n1482), .B1(n1680), .A0N(\gbuff[24][17] ), .A1N(n1681), 
        .Y(n2033) );
  OAI2BB2XL U1591 ( .B0(n1480), .B1(n1681), .A0N(\gbuff[24][18] ), .A1N(n1681), 
        .Y(n2032) );
  OAI2BB2XL U1592 ( .B0(n1478), .B1(n1680), .A0N(\gbuff[24][19] ), .A1N(n1681), 
        .Y(n2031) );
  OAI2BB2XL U1593 ( .B0(n1476), .B1(n1681), .A0N(\gbuff[24][20] ), .A1N(n1681), 
        .Y(n2030) );
  OAI2BB2XL U1594 ( .B0(n1474), .B1(n1680), .A0N(\gbuff[24][21] ), .A1N(n1681), 
        .Y(n2029) );
  OAI2BB2XL U1595 ( .B0(n1472), .B1(n1681), .A0N(\gbuff[24][22] ), .A1N(n1682), 
        .Y(n2028) );
  OAI2BB2XL U1596 ( .B0(n1470), .B1(n1681), .A0N(\gbuff[24][23] ), .A1N(n1681), 
        .Y(n2027) );
  OAI2BB2XL U1597 ( .B0(n1468), .B1(n1680), .A0N(\gbuff[24][24] ), .A1N(n1682), 
        .Y(n2026) );
  OAI2BB2XL U1598 ( .B0(n1466), .B1(n1681), .A0N(\gbuff[24][25] ), .A1N(n1682), 
        .Y(n2025) );
  OAI2BB2XL U1599 ( .B0(n1464), .B1(n1681), .A0N(\gbuff[24][26] ), .A1N(n1682), 
        .Y(n2024) );
  OAI2BB2XL U1600 ( .B0(n1462), .B1(n1681), .A0N(\gbuff[24][27] ), .A1N(n1682), 
        .Y(n2023) );
  OAI2BB2XL U1601 ( .B0(n1460), .B1(n1681), .A0N(\gbuff[24][28] ), .A1N(n1682), 
        .Y(n2022) );
  OAI2BB2XL U1602 ( .B0(n1458), .B1(n1681), .A0N(\gbuff[24][29] ), .A1N(n1682), 
        .Y(n2021) );
  OAI2BB2XL U1603 ( .B0(n1456), .B1(n1681), .A0N(\gbuff[24][30] ), .A1N(n1682), 
        .Y(n2020) );
  OAI2BB2XL U1604 ( .B0(n1454), .B1(n1681), .A0N(\gbuff[24][31] ), .A1N(n1680), 
        .Y(n2019) );
  OAI2BB2XL U1605 ( .B0(n1516), .B1(n1677), .A0N(\gbuff[25][0] ), .A1N(n1679), 
        .Y(n2018) );
  OAI2BB2XL U1606 ( .B0(n1514), .B1(n1677), .A0N(\gbuff[25][1] ), .A1N(n1678), 
        .Y(n2017) );
  OAI2BB2XL U1607 ( .B0(n1512), .B1(n1677), .A0N(\gbuff[25][2] ), .A1N(n1677), 
        .Y(n2016) );
  OAI2BB2XL U1608 ( .B0(n1510), .B1(n1677), .A0N(\gbuff[25][3] ), .A1N(n1679), 
        .Y(n2015) );
  OAI2BB2XL U1609 ( .B0(n1508), .B1(n1677), .A0N(\gbuff[25][4] ), .A1N(n1679), 
        .Y(n2014) );
  OAI2BB2XL U1610 ( .B0(n1506), .B1(n1677), .A0N(\gbuff[25][5] ), .A1N(n1679), 
        .Y(n2013) );
  OAI2BB2XL U1611 ( .B0(n1504), .B1(n1677), .A0N(\gbuff[25][6] ), .A1N(n1679), 
        .Y(n2012) );
  OAI2BB2XL U1612 ( .B0(n1502), .B1(n1677), .A0N(\gbuff[25][7] ), .A1N(n1679), 
        .Y(n2011) );
  OAI2BB2XL U1613 ( .B0(n1500), .B1(n1677), .A0N(\gbuff[25][8] ), .A1N(n1679), 
        .Y(n2010) );
  OAI2BB2XL U1614 ( .B0(n1498), .B1(n1677), .A0N(\gbuff[25][9] ), .A1N(n1679), 
        .Y(n2009) );
  OAI2BB2XL U1615 ( .B0(n1496), .B1(n1677), .A0N(\gbuff[25][10] ), .A1N(n1679), 
        .Y(n2008) );
  OAI2BB2XL U1616 ( .B0(n1494), .B1(n1677), .A0N(\gbuff[25][11] ), .A1N(n1679), 
        .Y(n2007) );
  OAI2BB2XL U1617 ( .B0(n1492), .B1(n1677), .A0N(\gbuff[25][12] ), .A1N(n1679), 
        .Y(n2006) );
  OAI2BB2XL U1618 ( .B0(n1490), .B1(n1677), .A0N(\gbuff[25][13] ), .A1N(n1679), 
        .Y(n2005) );
  OAI2BB2XL U1619 ( .B0(n1488), .B1(n1678), .A0N(\gbuff[25][14] ), .A1N(n1679), 
        .Y(n2004) );
  OAI2BB2XL U1620 ( .B0(n1486), .B1(n1677), .A0N(\gbuff[25][15] ), .A1N(n1678), 
        .Y(n2003) );
  OAI2BB2XL U1621 ( .B0(n1484), .B1(n1678), .A0N(\gbuff[25][16] ), .A1N(n1679), 
        .Y(n2002) );
  OAI2BB2XL U1622 ( .B0(n1482), .B1(n1677), .A0N(\gbuff[25][17] ), .A1N(n1678), 
        .Y(n2001) );
  OAI2BB2XL U1623 ( .B0(n1480), .B1(n1678), .A0N(\gbuff[25][18] ), .A1N(n1678), 
        .Y(n2000) );
  OAI2BB2XL U1624 ( .B0(n1478), .B1(n1677), .A0N(\gbuff[25][19] ), .A1N(n1678), 
        .Y(n1999) );
  OAI2BB2XL U1625 ( .B0(n1476), .B1(n1678), .A0N(\gbuff[25][20] ), .A1N(n1678), 
        .Y(n1998) );
  OAI2BB2XL U1626 ( .B0(n1474), .B1(n1677), .A0N(\gbuff[25][21] ), .A1N(n1678), 
        .Y(n1997) );
  OAI2BB2XL U1627 ( .B0(n1472), .B1(n1678), .A0N(\gbuff[25][22] ), .A1N(n1679), 
        .Y(n1996) );
  OAI2BB2XL U1628 ( .B0(n1470), .B1(n1678), .A0N(\gbuff[25][23] ), .A1N(n1678), 
        .Y(n1995) );
  OAI2BB2XL U1629 ( .B0(n1468), .B1(n1677), .A0N(\gbuff[25][24] ), .A1N(n1679), 
        .Y(n1994) );
  OAI2BB2XL U1630 ( .B0(n1466), .B1(n1678), .A0N(\gbuff[25][25] ), .A1N(n1679), 
        .Y(n1993) );
  OAI2BB2XL U1631 ( .B0(n1464), .B1(n1678), .A0N(\gbuff[25][26] ), .A1N(n1679), 
        .Y(n1992) );
  OAI2BB2XL U1632 ( .B0(n1462), .B1(n1678), .A0N(\gbuff[25][27] ), .A1N(n1679), 
        .Y(n1991) );
  OAI2BB2XL U1633 ( .B0(n1460), .B1(n1678), .A0N(\gbuff[25][28] ), .A1N(n1679), 
        .Y(n1990) );
  OAI2BB2XL U1634 ( .B0(n1458), .B1(n1678), .A0N(\gbuff[25][29] ), .A1N(n1679), 
        .Y(n1989) );
  OAI2BB2XL U1635 ( .B0(n1456), .B1(n1678), .A0N(\gbuff[25][30] ), .A1N(n1679), 
        .Y(n1988) );
  OAI2BB2XL U1636 ( .B0(n1454), .B1(n1678), .A0N(\gbuff[25][31] ), .A1N(n1677), 
        .Y(n1987) );
  OAI2BB2XL U1637 ( .B0(n1516), .B1(n1674), .A0N(\gbuff[26][0] ), .A1N(n1676), 
        .Y(n1986) );
  OAI2BB2XL U1638 ( .B0(n1514), .B1(n1674), .A0N(\gbuff[26][1] ), .A1N(n1675), 
        .Y(n1985) );
  OAI2BB2XL U1639 ( .B0(n1512), .B1(n1674), .A0N(\gbuff[26][2] ), .A1N(n1674), 
        .Y(n1984) );
  OAI2BB2XL U1640 ( .B0(n1510), .B1(n1674), .A0N(\gbuff[26][3] ), .A1N(n1676), 
        .Y(n1983) );
  OAI2BB2XL U1641 ( .B0(n1508), .B1(n1674), .A0N(\gbuff[26][4] ), .A1N(n1676), 
        .Y(n1982) );
  OAI2BB2XL U1642 ( .B0(n1506), .B1(n1674), .A0N(\gbuff[26][5] ), .A1N(n1676), 
        .Y(n1981) );
  OAI2BB2XL U1643 ( .B0(n1504), .B1(n1674), .A0N(\gbuff[26][6] ), .A1N(n1676), 
        .Y(n1980) );
  OAI2BB2XL U1644 ( .B0(n1502), .B1(n1674), .A0N(\gbuff[26][7] ), .A1N(n1676), 
        .Y(n1979) );
  OAI2BB2XL U1645 ( .B0(n1500), .B1(n1674), .A0N(\gbuff[26][8] ), .A1N(n1676), 
        .Y(n1978) );
  OAI2BB2XL U1646 ( .B0(n1498), .B1(n1674), .A0N(\gbuff[26][9] ), .A1N(n1676), 
        .Y(n1977) );
  OAI2BB2XL U1647 ( .B0(n1496), .B1(n1674), .A0N(\gbuff[26][10] ), .A1N(n1676), 
        .Y(n1976) );
  OAI2BB2XL U1648 ( .B0(n1494), .B1(n1674), .A0N(\gbuff[26][11] ), .A1N(n1676), 
        .Y(n1975) );
  OAI2BB2XL U1649 ( .B0(n1492), .B1(n1674), .A0N(\gbuff[26][12] ), .A1N(n1676), 
        .Y(n1974) );
  OAI2BB2XL U1650 ( .B0(n1490), .B1(n1674), .A0N(\gbuff[26][13] ), .A1N(n1676), 
        .Y(n1973) );
  OAI2BB2XL U1651 ( .B0(n1488), .B1(n1675), .A0N(\gbuff[26][14] ), .A1N(n1676), 
        .Y(n1972) );
  OAI2BB2XL U1652 ( .B0(n1486), .B1(n1674), .A0N(\gbuff[26][15] ), .A1N(n1675), 
        .Y(n1971) );
  OAI2BB2XL U1653 ( .B0(n1484), .B1(n1675), .A0N(\gbuff[26][16] ), .A1N(n1676), 
        .Y(n1970) );
  OAI2BB2XL U1654 ( .B0(n1482), .B1(n1674), .A0N(\gbuff[26][17] ), .A1N(n1675), 
        .Y(n1969) );
  OAI2BB2XL U1655 ( .B0(n1480), .B1(n1675), .A0N(\gbuff[26][18] ), .A1N(n1675), 
        .Y(n1968) );
  OAI2BB2XL U1656 ( .B0(n1478), .B1(n1674), .A0N(\gbuff[26][19] ), .A1N(n1675), 
        .Y(n1967) );
  OAI2BB2XL U1657 ( .B0(n1476), .B1(n1675), .A0N(\gbuff[26][20] ), .A1N(n1675), 
        .Y(n1966) );
  OAI2BB2XL U1658 ( .B0(n1474), .B1(n1674), .A0N(\gbuff[26][21] ), .A1N(n1675), 
        .Y(n1965) );
  OAI2BB2XL U1659 ( .B0(n1472), .B1(n1675), .A0N(\gbuff[26][22] ), .A1N(n1676), 
        .Y(n1964) );
  OAI2BB2XL U1660 ( .B0(n1470), .B1(n1675), .A0N(\gbuff[26][23] ), .A1N(n1675), 
        .Y(n1963) );
  OAI2BB2XL U1661 ( .B0(n1468), .B1(n1674), .A0N(\gbuff[26][24] ), .A1N(n1676), 
        .Y(n1962) );
  OAI2BB2XL U1662 ( .B0(n1466), .B1(n1675), .A0N(\gbuff[26][25] ), .A1N(n1676), 
        .Y(n1961) );
  OAI2BB2XL U1663 ( .B0(n1464), .B1(n1675), .A0N(\gbuff[26][26] ), .A1N(n1676), 
        .Y(n1960) );
  OAI2BB2XL U1664 ( .B0(n1462), .B1(n1675), .A0N(\gbuff[26][27] ), .A1N(n1676), 
        .Y(n1959) );
  OAI2BB2XL U1665 ( .B0(n1460), .B1(n1675), .A0N(\gbuff[26][28] ), .A1N(n1676), 
        .Y(n1958) );
  OAI2BB2XL U1666 ( .B0(n1458), .B1(n1675), .A0N(\gbuff[26][29] ), .A1N(n1676), 
        .Y(n1957) );
  OAI2BB2XL U1667 ( .B0(n1456), .B1(n1675), .A0N(\gbuff[26][30] ), .A1N(n1676), 
        .Y(n1956) );
  OAI2BB2XL U1668 ( .B0(n1454), .B1(n1675), .A0N(\gbuff[26][31] ), .A1N(n1674), 
        .Y(n1955) );
  OAI2BB2XL U1669 ( .B0(n1516), .B1(n1671), .A0N(\gbuff[27][0] ), .A1N(n1673), 
        .Y(n1954) );
  OAI2BB2XL U1670 ( .B0(n1514), .B1(n1671), .A0N(\gbuff[27][1] ), .A1N(n1672), 
        .Y(n1953) );
  OAI2BB2XL U1671 ( .B0(n1512), .B1(n1671), .A0N(\gbuff[27][2] ), .A1N(n1671), 
        .Y(n1952) );
  OAI2BB2XL U1672 ( .B0(n1510), .B1(n1671), .A0N(\gbuff[27][3] ), .A1N(n1673), 
        .Y(n1951) );
  OAI2BB2XL U1673 ( .B0(n1508), .B1(n1671), .A0N(\gbuff[27][4] ), .A1N(n1673), 
        .Y(n1950) );
  OAI2BB2XL U1674 ( .B0(n1506), .B1(n1671), .A0N(\gbuff[27][5] ), .A1N(n1673), 
        .Y(n1949) );
  OAI2BB2XL U1675 ( .B0(n1504), .B1(n1671), .A0N(\gbuff[27][6] ), .A1N(n1673), 
        .Y(n1948) );
  OAI2BB2XL U1676 ( .B0(n1502), .B1(n1671), .A0N(\gbuff[27][7] ), .A1N(n1673), 
        .Y(n1947) );
  OAI2BB2XL U1677 ( .B0(n1500), .B1(n1671), .A0N(\gbuff[27][8] ), .A1N(n1673), 
        .Y(n1946) );
  OAI2BB2XL U1678 ( .B0(n1498), .B1(n1671), .A0N(\gbuff[27][9] ), .A1N(n1673), 
        .Y(n1945) );
  OAI2BB2XL U1679 ( .B0(n1496), .B1(n1671), .A0N(\gbuff[27][10] ), .A1N(n1673), 
        .Y(n1944) );
  OAI2BB2XL U1680 ( .B0(n1494), .B1(n1671), .A0N(\gbuff[27][11] ), .A1N(n1673), 
        .Y(n1943) );
  OAI2BB2XL U1681 ( .B0(n1492), .B1(n1671), .A0N(\gbuff[27][12] ), .A1N(n1673), 
        .Y(n1942) );
  OAI2BB2XL U1682 ( .B0(n1490), .B1(n1671), .A0N(\gbuff[27][13] ), .A1N(n1673), 
        .Y(n1941) );
  OAI2BB2XL U1683 ( .B0(n1488), .B1(n1672), .A0N(\gbuff[27][14] ), .A1N(n1673), 
        .Y(n1940) );
  OAI2BB2XL U1684 ( .B0(n1486), .B1(n1671), .A0N(\gbuff[27][15] ), .A1N(n1672), 
        .Y(n1939) );
  OAI2BB2XL U1685 ( .B0(n1484), .B1(n1672), .A0N(\gbuff[27][16] ), .A1N(n1673), 
        .Y(n1938) );
  OAI2BB2XL U1686 ( .B0(n1482), .B1(n1671), .A0N(\gbuff[27][17] ), .A1N(n1672), 
        .Y(n1937) );
  OAI2BB2XL U1687 ( .B0(n1480), .B1(n1672), .A0N(\gbuff[27][18] ), .A1N(n1672), 
        .Y(n1936) );
  OAI2BB2XL U1688 ( .B0(n1478), .B1(n1671), .A0N(\gbuff[27][19] ), .A1N(n1672), 
        .Y(n1935) );
  OAI2BB2XL U1689 ( .B0(n1476), .B1(n1672), .A0N(\gbuff[27][20] ), .A1N(n1672), 
        .Y(n1934) );
  OAI2BB2XL U1690 ( .B0(n1474), .B1(n1671), .A0N(\gbuff[27][21] ), .A1N(n1672), 
        .Y(n1933) );
  OAI2BB2XL U1691 ( .B0(n1472), .B1(n1672), .A0N(\gbuff[27][22] ), .A1N(n1673), 
        .Y(n1932) );
  OAI2BB2XL U1692 ( .B0(n1470), .B1(n1672), .A0N(\gbuff[27][23] ), .A1N(n1672), 
        .Y(n1931) );
  OAI2BB2XL U1693 ( .B0(n1468), .B1(n1671), .A0N(\gbuff[27][24] ), .A1N(n1673), 
        .Y(n1930) );
  OAI2BB2XL U1694 ( .B0(n1466), .B1(n1672), .A0N(\gbuff[27][25] ), .A1N(n1673), 
        .Y(n1929) );
  OAI2BB2XL U1695 ( .B0(n1464), .B1(n1672), .A0N(\gbuff[27][26] ), .A1N(n1673), 
        .Y(n1928) );
  OAI2BB2XL U1696 ( .B0(n1462), .B1(n1672), .A0N(\gbuff[27][27] ), .A1N(n1673), 
        .Y(n1927) );
  OAI2BB2XL U1697 ( .B0(n1460), .B1(n1672), .A0N(\gbuff[27][28] ), .A1N(n1673), 
        .Y(n1926) );
  OAI2BB2XL U1698 ( .B0(n1458), .B1(n1672), .A0N(\gbuff[27][29] ), .A1N(n1673), 
        .Y(n1925) );
  OAI2BB2XL U1699 ( .B0(n1456), .B1(n1672), .A0N(\gbuff[27][30] ), .A1N(n1673), 
        .Y(n1924) );
  OAI2BB2XL U1700 ( .B0(n1454), .B1(n1672), .A0N(\gbuff[27][31] ), .A1N(n1671), 
        .Y(n1923) );
  OAI2BB2XL U1701 ( .B0(n1516), .B1(n1668), .A0N(\gbuff[28][0] ), .A1N(n1669), 
        .Y(n1922) );
  OAI2BB2XL U1702 ( .B0(n1514), .B1(n1668), .A0N(\gbuff[28][1] ), .A1N(n1668), 
        .Y(n1921) );
  OAI2BB2XL U1703 ( .B0(n1512), .B1(n1668), .A0N(\gbuff[28][2] ), .A1N(n1670), 
        .Y(n1920) );
  OAI2BB2XL U1704 ( .B0(n1510), .B1(n1668), .A0N(\gbuff[28][3] ), .A1N(n1670), 
        .Y(n1919) );
  OAI2BB2XL U1705 ( .B0(n1508), .B1(n1668), .A0N(\gbuff[28][4] ), .A1N(n1668), 
        .Y(n1918) );
  OAI2BB2XL U1706 ( .B0(n1506), .B1(n1668), .A0N(\gbuff[28][5] ), .A1N(n1670), 
        .Y(n1917) );
  OAI2BB2XL U1707 ( .B0(n1504), .B1(n1668), .A0N(\gbuff[28][6] ), .A1N(n1670), 
        .Y(n1916) );
  OAI2BB2XL U1708 ( .B0(n1502), .B1(n1668), .A0N(\gbuff[28][7] ), .A1N(n1670), 
        .Y(n1915) );
  OAI2BB2XL U1709 ( .B0(n1500), .B1(n1668), .A0N(\gbuff[28][8] ), .A1N(n1670), 
        .Y(n1914) );
  OAI2BB2XL U1710 ( .B0(n1498), .B1(n1668), .A0N(\gbuff[28][9] ), .A1N(n1670), 
        .Y(n1913) );
  OAI2BB2XL U1711 ( .B0(n1496), .B1(n1668), .A0N(\gbuff[28][10] ), .A1N(n1670), 
        .Y(n1912) );
  OAI2BB2XL U1712 ( .B0(n1494), .B1(n1668), .A0N(\gbuff[28][11] ), .A1N(n1670), 
        .Y(n1911) );
  OAI2BB2XL U1713 ( .B0(n1492), .B1(n1668), .A0N(\gbuff[28][12] ), .A1N(n1670), 
        .Y(n1910) );
  OAI2BB2XL U1714 ( .B0(n1490), .B1(n1668), .A0N(\gbuff[28][13] ), .A1N(n1670), 
        .Y(n1909) );
  OAI2BB2XL U1715 ( .B0(n1488), .B1(n1668), .A0N(\gbuff[28][14] ), .A1N(n1670), 
        .Y(n1908) );
  OAI2BB2XL U1716 ( .B0(n1486), .B1(n1668), .A0N(\gbuff[28][15] ), .A1N(n1669), 
        .Y(n1907) );
  OAI2BB2XL U1717 ( .B0(n1484), .B1(n1668), .A0N(\gbuff[28][16] ), .A1N(n1670), 
        .Y(n1906) );
  OAI2BB2XL U1718 ( .B0(n1482), .B1(n1669), .A0N(\gbuff[28][17] ), .A1N(n1669), 
        .Y(n1905) );
  OAI2BB2XL U1719 ( .B0(n1480), .B1(n1668), .A0N(\gbuff[28][18] ), .A1N(n1669), 
        .Y(n1904) );
  OAI2BB2XL U1720 ( .B0(n1478), .B1(n1669), .A0N(\gbuff[28][19] ), .A1N(n1669), 
        .Y(n1903) );
  OAI2BB2XL U1721 ( .B0(n1476), .B1(n1668), .A0N(\gbuff[28][20] ), .A1N(n1669), 
        .Y(n1902) );
  OAI2BB2XL U1722 ( .B0(n1474), .B1(n1669), .A0N(\gbuff[28][21] ), .A1N(n1669), 
        .Y(n1901) );
  OAI2BB2XL U1723 ( .B0(n1472), .B1(n1669), .A0N(\gbuff[28][22] ), .A1N(n1670), 
        .Y(n1900) );
  OAI2BB2XL U1724 ( .B0(n1470), .B1(n1669), .A0N(\gbuff[28][23] ), .A1N(n1669), 
        .Y(n1899) );
  OAI2BB2XL U1725 ( .B0(n1468), .B1(n1670), .A0N(\gbuff[28][24] ), .A1N(n1670), 
        .Y(n1898) );
  OAI2BB2XL U1726 ( .B0(n1466), .B1(n1669), .A0N(\gbuff[28][25] ), .A1N(n1670), 
        .Y(n1897) );
  OAI2BB2XL U1727 ( .B0(n1464), .B1(n1669), .A0N(\gbuff[28][26] ), .A1N(n1670), 
        .Y(n1896) );
  OAI2BB2XL U1728 ( .B0(n1462), .B1(n1669), .A0N(\gbuff[28][27] ), .A1N(n1670), 
        .Y(n1895) );
  OAI2BB2XL U1729 ( .B0(n1460), .B1(n1669), .A0N(\gbuff[28][28] ), .A1N(n1670), 
        .Y(n1894) );
  OAI2BB2XL U1730 ( .B0(n1458), .B1(n1669), .A0N(\gbuff[28][29] ), .A1N(n1670), 
        .Y(n1893) );
  OAI2BB2XL U1731 ( .B0(n1456), .B1(n1669), .A0N(\gbuff[28][30] ), .A1N(n2822), 
        .Y(n1892) );
  OAI2BB2XL U1732 ( .B0(n1454), .B1(n1669), .A0N(\gbuff[28][31] ), .A1N(n2822), 
        .Y(n1891) );
  OAI2BB2XL U1733 ( .B0(n1516), .B1(n1665), .A0N(\gbuff[29][0] ), .A1N(n1667), 
        .Y(n1890) );
  OAI2BB2XL U1734 ( .B0(n1514), .B1(n1665), .A0N(\gbuff[29][1] ), .A1N(n2821), 
        .Y(n1889) );
  OAI2BB2XL U1735 ( .B0(n1512), .B1(n1665), .A0N(\gbuff[29][2] ), .A1N(n1665), 
        .Y(n1888) );
  OAI2BB2XL U1736 ( .B0(n1510), .B1(n1665), .A0N(\gbuff[29][3] ), .A1N(n1667), 
        .Y(n1887) );
  OAI2BB2XL U1737 ( .B0(n1508), .B1(n1665), .A0N(\gbuff[29][4] ), .A1N(n1667), 
        .Y(n1886) );
  OAI2BB2XL U1738 ( .B0(n1506), .B1(n1665), .A0N(\gbuff[29][5] ), .A1N(n1667), 
        .Y(n1885) );
  OAI2BB2XL U1739 ( .B0(n1504), .B1(n1665), .A0N(\gbuff[29][6] ), .A1N(n1667), 
        .Y(n1884) );
  OAI2BB2XL U1740 ( .B0(n1502), .B1(n1665), .A0N(\gbuff[29][7] ), .A1N(n1667), 
        .Y(n1883) );
  OAI2BB2XL U1741 ( .B0(n1500), .B1(n1665), .A0N(\gbuff[29][8] ), .A1N(n1667), 
        .Y(n1882) );
  OAI2BB2XL U1742 ( .B0(n1498), .B1(n1665), .A0N(\gbuff[29][9] ), .A1N(n1667), 
        .Y(n1881) );
  OAI2BB2XL U1743 ( .B0(n1496), .B1(n1665), .A0N(\gbuff[29][10] ), .A1N(n1667), 
        .Y(n1880) );
  OAI2BB2XL U1744 ( .B0(n1494), .B1(n1665), .A0N(\gbuff[29][11] ), .A1N(n1667), 
        .Y(n1879) );
  OAI2BB2XL U1745 ( .B0(n1492), .B1(n1665), .A0N(\gbuff[29][12] ), .A1N(n1667), 
        .Y(n1878) );
  OAI2BB2XL U1746 ( .B0(n1490), .B1(n1665), .A0N(\gbuff[29][13] ), .A1N(n1667), 
        .Y(n1877) );
  OAI2BB2XL U1747 ( .B0(n1488), .B1(n1666), .A0N(\gbuff[29][14] ), .A1N(n1667), 
        .Y(n1876) );
  OAI2BB2XL U1748 ( .B0(n1486), .B1(n1665), .A0N(\gbuff[29][15] ), .A1N(n1666), 
        .Y(n1875) );
  OAI2BB2XL U1749 ( .B0(n1484), .B1(n1666), .A0N(\gbuff[29][16] ), .A1N(n1667), 
        .Y(n1874) );
  OAI2BB2XL U1750 ( .B0(n1482), .B1(n1665), .A0N(\gbuff[29][17] ), .A1N(n1666), 
        .Y(n1873) );
  OAI2BB2XL U1751 ( .B0(n1480), .B1(n1666), .A0N(\gbuff[29][18] ), .A1N(n1666), 
        .Y(n1872) );
  OAI2BB2XL U1752 ( .B0(n1478), .B1(n1665), .A0N(\gbuff[29][19] ), .A1N(n1666), 
        .Y(n1871) );
  OAI2BB2XL U1753 ( .B0(n1476), .B1(n1666), .A0N(\gbuff[29][20] ), .A1N(n1666), 
        .Y(n1870) );
  OAI2BB2XL U1754 ( .B0(n1474), .B1(n1665), .A0N(\gbuff[29][21] ), .A1N(n1666), 
        .Y(n1869) );
  OAI2BB2XL U1755 ( .B0(n1472), .B1(n1666), .A0N(\gbuff[29][22] ), .A1N(n1667), 
        .Y(n1868) );
  OAI2BB2XL U1756 ( .B0(n1470), .B1(n1666), .A0N(\gbuff[29][23] ), .A1N(n1666), 
        .Y(n1867) );
  OAI2BB2XL U1757 ( .B0(n1468), .B1(n2821), .A0N(\gbuff[29][24] ), .A1N(n1667), 
        .Y(n1866) );
  OAI2BB2XL U1758 ( .B0(n1466), .B1(n1666), .A0N(\gbuff[29][25] ), .A1N(n1667), 
        .Y(n1865) );
  OAI2BB2XL U1759 ( .B0(n1464), .B1(n1666), .A0N(\gbuff[29][26] ), .A1N(n1667), 
        .Y(n1864) );
  OAI2BB2XL U1760 ( .B0(n1462), .B1(n1666), .A0N(\gbuff[29][27] ), .A1N(n1667), 
        .Y(n1863) );
  OAI2BB2XL U1761 ( .B0(n1460), .B1(n1666), .A0N(\gbuff[29][28] ), .A1N(n1667), 
        .Y(n1862) );
  OAI2BB2XL U1762 ( .B0(n1458), .B1(n1666), .A0N(\gbuff[29][29] ), .A1N(n1667), 
        .Y(n1861) );
  OAI2BB2XL U1763 ( .B0(n1456), .B1(n1666), .A0N(\gbuff[29][30] ), .A1N(n1667), 
        .Y(n1860) );
  OAI2BB2XL U1764 ( .B0(n1454), .B1(n1666), .A0N(\gbuff[29][31] ), .A1N(n1665), 
        .Y(n1859) );
  OAI2BB2XL U1765 ( .B0(n1516), .B1(n1662), .A0N(\gbuff[30][0] ), .A1N(n1664), 
        .Y(n1858) );
  OAI2BB2XL U1766 ( .B0(n1514), .B1(n1662), .A0N(\gbuff[30][1] ), .A1N(n2820), 
        .Y(n1857) );
  OAI2BB2XL U1767 ( .B0(n1512), .B1(n1662), .A0N(\gbuff[30][2] ), .A1N(n1662), 
        .Y(n1856) );
  OAI2BB2XL U1768 ( .B0(n1510), .B1(n1662), .A0N(\gbuff[30][3] ), .A1N(n1664), 
        .Y(n1855) );
  OAI2BB2XL U1769 ( .B0(n1508), .B1(n1662), .A0N(\gbuff[30][4] ), .A1N(n1664), 
        .Y(n1854) );
  OAI2BB2XL U1770 ( .B0(n1506), .B1(n1662), .A0N(\gbuff[30][5] ), .A1N(n1664), 
        .Y(n1853) );
  OAI2BB2XL U1771 ( .B0(n1504), .B1(n1662), .A0N(\gbuff[30][6] ), .A1N(n1664), 
        .Y(n1852) );
  OAI2BB2XL U1772 ( .B0(n1502), .B1(n1662), .A0N(\gbuff[30][7] ), .A1N(n1664), 
        .Y(n1851) );
  OAI2BB2XL U1773 ( .B0(n1500), .B1(n1662), .A0N(\gbuff[30][8] ), .A1N(n1664), 
        .Y(n1850) );
  OAI2BB2XL U1774 ( .B0(n1498), .B1(n1662), .A0N(\gbuff[30][9] ), .A1N(n1664), 
        .Y(n1849) );
  OAI2BB2XL U1775 ( .B0(n1496), .B1(n1662), .A0N(\gbuff[30][10] ), .A1N(n1664), 
        .Y(n1848) );
  OAI2BB2XL U1776 ( .B0(n1494), .B1(n1662), .A0N(\gbuff[30][11] ), .A1N(n1664), 
        .Y(n1847) );
  OAI2BB2XL U1777 ( .B0(n1492), .B1(n1662), .A0N(\gbuff[30][12] ), .A1N(n1664), 
        .Y(n1846) );
  OAI2BB2XL U1778 ( .B0(n1490), .B1(n1662), .A0N(\gbuff[30][13] ), .A1N(n1664), 
        .Y(n1845) );
  OAI2BB2XL U1779 ( .B0(n1488), .B1(n1663), .A0N(\gbuff[30][14] ), .A1N(n1664), 
        .Y(n1844) );
  OAI2BB2XL U1780 ( .B0(n1486), .B1(n1662), .A0N(\gbuff[30][15] ), .A1N(n1663), 
        .Y(n1843) );
  OAI2BB2XL U1781 ( .B0(n1484), .B1(n1663), .A0N(\gbuff[30][16] ), .A1N(n1664), 
        .Y(n1842) );
  OAI2BB2XL U1782 ( .B0(n1482), .B1(n1662), .A0N(\gbuff[30][17] ), .A1N(n1663), 
        .Y(n1841) );
  OAI2BB2XL U1783 ( .B0(n1480), .B1(n1663), .A0N(\gbuff[30][18] ), .A1N(n1663), 
        .Y(n1840) );
  OAI2BB2XL U1784 ( .B0(n1478), .B1(n1662), .A0N(\gbuff[30][19] ), .A1N(n1663), 
        .Y(n1839) );
  OAI2BB2XL U1785 ( .B0(n1476), .B1(n1663), .A0N(\gbuff[30][20] ), .A1N(n1663), 
        .Y(n1838) );
  OAI2BB2XL U1786 ( .B0(n1474), .B1(n1662), .A0N(\gbuff[30][21] ), .A1N(n1663), 
        .Y(n1837) );
  OAI2BB2XL U1787 ( .B0(n1472), .B1(n1663), .A0N(\gbuff[30][22] ), .A1N(n1664), 
        .Y(n1836) );
  OAI2BB2XL U1788 ( .B0(n1470), .B1(n1663), .A0N(\gbuff[30][23] ), .A1N(n1663), 
        .Y(n1835) );
  OAI2BB2XL U1789 ( .B0(n1468), .B1(n2820), .A0N(\gbuff[30][24] ), .A1N(n1664), 
        .Y(n1834) );
  OAI2BB2XL U1790 ( .B0(n1466), .B1(n1663), .A0N(\gbuff[30][25] ), .A1N(n1664), 
        .Y(n1833) );
  OAI2BB2XL U1791 ( .B0(n1464), .B1(n1663), .A0N(\gbuff[30][26] ), .A1N(n1664), 
        .Y(n1832) );
  OAI2BB2XL U1792 ( .B0(n1462), .B1(n1663), .A0N(\gbuff[30][27] ), .A1N(n1664), 
        .Y(n1831) );
  OAI2BB2XL U1793 ( .B0(n1460), .B1(n1663), .A0N(\gbuff[30][28] ), .A1N(n1664), 
        .Y(n1830) );
  OAI2BB2XL U1794 ( .B0(n1458), .B1(n1663), .A0N(\gbuff[30][29] ), .A1N(n1664), 
        .Y(n1829) );
  OAI2BB2XL U1795 ( .B0(n1456), .B1(n1663), .A0N(\gbuff[30][30] ), .A1N(n1664), 
        .Y(n1828) );
  OAI2BB2XL U1796 ( .B0(n1454), .B1(n1663), .A0N(\gbuff[30][31] ), .A1N(n1662), 
        .Y(n1827) );
  OAI2BB2XL U1797 ( .B0(n1516), .B1(n1659), .A0N(\gbuff[31][0] ), .A1N(n1661), 
        .Y(n1826) );
  OAI2BB2XL U1798 ( .B0(n1514), .B1(n1659), .A0N(\gbuff[31][1] ), .A1N(n2819), 
        .Y(n1825) );
  OAI2BB2XL U1799 ( .B0(n1512), .B1(n1659), .A0N(\gbuff[31][2] ), .A1N(n1659), 
        .Y(n1824) );
  OAI2BB2XL U1800 ( .B0(n1510), .B1(n1659), .A0N(\gbuff[31][3] ), .A1N(n1661), 
        .Y(n1823) );
  OAI2BB2XL U1801 ( .B0(n1508), .B1(n1659), .A0N(\gbuff[31][4] ), .A1N(n1661), 
        .Y(n1822) );
  OAI2BB2XL U1802 ( .B0(n1506), .B1(n1659), .A0N(\gbuff[31][5] ), .A1N(n1661), 
        .Y(n1821) );
  OAI2BB2XL U1803 ( .B0(n1504), .B1(n1659), .A0N(\gbuff[31][6] ), .A1N(n1661), 
        .Y(n1820) );
  OAI2BB2XL U1804 ( .B0(n1502), .B1(n1659), .A0N(\gbuff[31][7] ), .A1N(n1661), 
        .Y(n1819) );
  OAI2BB2XL U1805 ( .B0(n1500), .B1(n1659), .A0N(\gbuff[31][8] ), .A1N(n1661), 
        .Y(n1818) );
  OAI2BB2XL U1806 ( .B0(n1498), .B1(n1659), .A0N(\gbuff[31][9] ), .A1N(n1661), 
        .Y(n1817) );
  OAI2BB2XL U1807 ( .B0(n1496), .B1(n1659), .A0N(\gbuff[31][10] ), .A1N(n1661), 
        .Y(n1816) );
  OAI2BB2XL U1808 ( .B0(n1494), .B1(n1659), .A0N(\gbuff[31][11] ), .A1N(n1661), 
        .Y(n1815) );
  OAI2BB2XL U1809 ( .B0(n1492), .B1(n1659), .A0N(\gbuff[31][12] ), .A1N(n1661), 
        .Y(n1814) );
  OAI2BB2XL U1810 ( .B0(n1490), .B1(n1659), .A0N(\gbuff[31][13] ), .A1N(n1661), 
        .Y(n1813) );
  OAI2BB2XL U1811 ( .B0(n1488), .B1(n1660), .A0N(\gbuff[31][14] ), .A1N(n1661), 
        .Y(n1812) );
  OAI2BB2XL U1812 ( .B0(n1486), .B1(n1659), .A0N(\gbuff[31][15] ), .A1N(n1660), 
        .Y(n1811) );
  OAI2BB2XL U1813 ( .B0(n1484), .B1(n1660), .A0N(\gbuff[31][16] ), .A1N(n1661), 
        .Y(n1810) );
  OAI2BB2XL U1814 ( .B0(n1482), .B1(n1659), .A0N(\gbuff[31][17] ), .A1N(n1660), 
        .Y(n1809) );
  OAI2BB2XL U1815 ( .B0(n1480), .B1(n1660), .A0N(\gbuff[31][18] ), .A1N(n1660), 
        .Y(n1808) );
  OAI2BB2XL U1816 ( .B0(n1478), .B1(n1659), .A0N(\gbuff[31][19] ), .A1N(n1660), 
        .Y(n1807) );
  OAI2BB2XL U1817 ( .B0(n1476), .B1(n1660), .A0N(\gbuff[31][20] ), .A1N(n1660), 
        .Y(n1806) );
  OAI2BB2XL U1818 ( .B0(n1474), .B1(n1659), .A0N(\gbuff[31][21] ), .A1N(n1660), 
        .Y(n1805) );
  OAI2BB2XL U1819 ( .B0(n1472), .B1(n1660), .A0N(\gbuff[31][22] ), .A1N(n1661), 
        .Y(n1804) );
  OAI2BB2XL U1820 ( .B0(n1470), .B1(n1660), .A0N(\gbuff[31][23] ), .A1N(n1660), 
        .Y(n1803) );
  OAI2BB2XL U1821 ( .B0(n1468), .B1(n2819), .A0N(\gbuff[31][24] ), .A1N(n1661), 
        .Y(n1802) );
  OAI2BB2XL U1822 ( .B0(n1466), .B1(n1660), .A0N(\gbuff[31][25] ), .A1N(n1661), 
        .Y(n1801) );
  OAI2BB2XL U1823 ( .B0(n1464), .B1(n1660), .A0N(\gbuff[31][26] ), .A1N(n1661), 
        .Y(n1800) );
  OAI2BB2XL U1824 ( .B0(n1462), .B1(n1660), .A0N(\gbuff[31][27] ), .A1N(n1661), 
        .Y(n1799) );
  OAI2BB2XL U1825 ( .B0(n1460), .B1(n1660), .A0N(\gbuff[31][28] ), .A1N(n1661), 
        .Y(n1798) );
  OAI2BB2XL U1826 ( .B0(n1458), .B1(n1660), .A0N(\gbuff[31][29] ), .A1N(n1661), 
        .Y(n1797) );
  OAI2BB2XL U1827 ( .B0(n1456), .B1(n1660), .A0N(\gbuff[31][30] ), .A1N(n1661), 
        .Y(n1796) );
  OAI2BB2XL U1828 ( .B0(n1454), .B1(n1660), .A0N(\gbuff[31][31] ), .A1N(n1659), 
        .Y(n1795) );
endmodule


module global_buffer_1 ( clk, rst, wr_en, index, data_in, data_out );
  input [7:0] index;
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, wr_en;
  wire   N10, N11, N12, N13, N14, \gbuff[1][31] , \gbuff[1][30] ,
         \gbuff[1][29] , \gbuff[1][28] , \gbuff[1][27] , \gbuff[1][26] ,
         \gbuff[1][25] , \gbuff[1][24] , \gbuff[1][23] , \gbuff[1][22] ,
         \gbuff[1][21] , \gbuff[1][20] , \gbuff[1][19] , \gbuff[1][18] ,
         \gbuff[1][17] , \gbuff[1][16] , \gbuff[1][15] , \gbuff[1][14] ,
         \gbuff[1][13] , \gbuff[1][12] , \gbuff[1][11] , \gbuff[1][10] ,
         \gbuff[1][9] , \gbuff[1][8] , \gbuff[1][7] , \gbuff[1][6] ,
         \gbuff[1][5] , \gbuff[1][4] , \gbuff[1][3] , \gbuff[1][2] ,
         \gbuff[1][1] , \gbuff[1][0] , \gbuff[0][31] , \gbuff[0][30] ,
         \gbuff[0][29] , \gbuff[0][28] , \gbuff[0][27] , \gbuff[0][26] ,
         \gbuff[0][25] , \gbuff[0][24] , \gbuff[0][23] , \gbuff[0][22] ,
         \gbuff[0][21] , \gbuff[0][20] , \gbuff[0][19] , \gbuff[0][18] ,
         \gbuff[0][17] , \gbuff[0][16] , \gbuff[0][15] , \gbuff[0][14] ,
         \gbuff[0][13] , \gbuff[0][12] , \gbuff[0][11] , \gbuff[0][10] ,
         \gbuff[0][9] , \gbuff[0][8] , \gbuff[0][7] , \gbuff[0][6] ,
         \gbuff[0][5] , \gbuff[0][4] , \gbuff[0][3] , \gbuff[0][2] ,
         \gbuff[0][1] , \gbuff[0][0] , \gbuff[3][31] , \gbuff[3][30] ,
         \gbuff[3][29] , \gbuff[3][28] , \gbuff[3][27] , \gbuff[3][26] ,
         \gbuff[3][25] , \gbuff[3][24] , \gbuff[3][23] , \gbuff[3][22] ,
         \gbuff[3][21] , \gbuff[3][20] , \gbuff[3][19] , \gbuff[3][18] ,
         \gbuff[3][17] , \gbuff[3][16] , \gbuff[3][15] , \gbuff[3][14] ,
         \gbuff[3][13] , \gbuff[3][12] , \gbuff[3][11] , \gbuff[3][10] ,
         \gbuff[3][9] , \gbuff[3][8] , \gbuff[3][7] , \gbuff[3][6] ,
         \gbuff[3][5] , \gbuff[3][4] , \gbuff[3][3] , \gbuff[3][2] ,
         \gbuff[3][1] , \gbuff[3][0] , \gbuff[2][31] , \gbuff[2][30] ,
         \gbuff[2][29] , \gbuff[2][28] , \gbuff[2][27] , \gbuff[2][26] ,
         \gbuff[2][25] , \gbuff[2][24] , \gbuff[2][23] , \gbuff[2][22] ,
         \gbuff[2][21] , \gbuff[2][20] , \gbuff[2][19] , \gbuff[2][18] ,
         \gbuff[2][17] , \gbuff[2][16] , \gbuff[2][15] , \gbuff[2][14] ,
         \gbuff[2][13] , \gbuff[2][12] , \gbuff[2][11] , \gbuff[2][10] ,
         \gbuff[2][9] , \gbuff[2][8] , \gbuff[2][7] , \gbuff[2][6] ,
         \gbuff[2][5] , \gbuff[2][4] , \gbuff[2][3] , \gbuff[2][2] ,
         \gbuff[2][1] , \gbuff[2][0] , \gbuff[5][31] , \gbuff[5][30] ,
         \gbuff[5][29] , \gbuff[5][28] , \gbuff[5][27] , \gbuff[5][26] ,
         \gbuff[5][25] , \gbuff[5][24] , \gbuff[5][23] , \gbuff[5][22] ,
         \gbuff[5][21] , \gbuff[5][20] , \gbuff[5][19] , \gbuff[5][18] ,
         \gbuff[5][17] , \gbuff[5][16] , \gbuff[5][15] , \gbuff[5][14] ,
         \gbuff[5][13] , \gbuff[5][12] , \gbuff[5][11] , \gbuff[5][10] ,
         \gbuff[5][9] , \gbuff[5][8] , \gbuff[5][7] , \gbuff[5][6] ,
         \gbuff[5][5] , \gbuff[5][4] , \gbuff[5][3] , \gbuff[5][2] ,
         \gbuff[5][1] , \gbuff[5][0] , \gbuff[4][31] , \gbuff[4][30] ,
         \gbuff[4][29] , \gbuff[4][28] , \gbuff[4][27] , \gbuff[4][26] ,
         \gbuff[4][25] , \gbuff[4][24] , \gbuff[4][23] , \gbuff[4][22] ,
         \gbuff[4][21] , \gbuff[4][20] , \gbuff[4][19] , \gbuff[4][18] ,
         \gbuff[4][17] , \gbuff[4][16] , \gbuff[4][15] , \gbuff[4][14] ,
         \gbuff[4][13] , \gbuff[4][12] , \gbuff[4][11] , \gbuff[4][10] ,
         \gbuff[4][9] , \gbuff[4][8] , \gbuff[4][7] , \gbuff[4][6] ,
         \gbuff[4][5] , \gbuff[4][4] , \gbuff[4][3] , \gbuff[4][2] ,
         \gbuff[4][1] , \gbuff[4][0] , \gbuff[7][31] , \gbuff[7][30] ,
         \gbuff[7][29] , \gbuff[7][28] , \gbuff[7][27] , \gbuff[7][26] ,
         \gbuff[7][25] , \gbuff[7][24] , \gbuff[7][23] , \gbuff[7][22] ,
         \gbuff[7][21] , \gbuff[7][20] , \gbuff[7][19] , \gbuff[7][18] ,
         \gbuff[7][17] , \gbuff[7][16] , \gbuff[7][15] , \gbuff[7][14] ,
         \gbuff[7][13] , \gbuff[7][12] , \gbuff[7][11] , \gbuff[7][10] ,
         \gbuff[7][9] , \gbuff[7][8] , \gbuff[7][7] , \gbuff[7][6] ,
         \gbuff[7][5] , \gbuff[7][4] , \gbuff[7][3] , \gbuff[7][2] ,
         \gbuff[7][1] , \gbuff[7][0] , \gbuff[6][31] , \gbuff[6][30] ,
         \gbuff[6][29] , \gbuff[6][28] , \gbuff[6][27] , \gbuff[6][26] ,
         \gbuff[6][25] , \gbuff[6][24] , \gbuff[6][23] , \gbuff[6][22] ,
         \gbuff[6][21] , \gbuff[6][20] , \gbuff[6][19] , \gbuff[6][18] ,
         \gbuff[6][17] , \gbuff[6][16] , \gbuff[6][15] , \gbuff[6][14] ,
         \gbuff[6][13] , \gbuff[6][12] , \gbuff[6][11] , \gbuff[6][10] ,
         \gbuff[6][9] , \gbuff[6][8] , \gbuff[6][7] , \gbuff[6][6] ,
         \gbuff[6][5] , \gbuff[6][4] , \gbuff[6][3] , \gbuff[6][2] ,
         \gbuff[6][1] , \gbuff[6][0] , \gbuff[9][31] , \gbuff[9][30] ,
         \gbuff[9][29] , \gbuff[9][28] , \gbuff[9][27] , \gbuff[9][26] ,
         \gbuff[9][25] , \gbuff[9][24] , \gbuff[9][23] , \gbuff[9][22] ,
         \gbuff[9][21] , \gbuff[9][20] , \gbuff[9][19] , \gbuff[9][18] ,
         \gbuff[9][17] , \gbuff[9][16] , \gbuff[9][15] , \gbuff[9][14] ,
         \gbuff[9][13] , \gbuff[9][12] , \gbuff[9][11] , \gbuff[9][10] ,
         \gbuff[9][9] , \gbuff[9][8] , \gbuff[9][7] , \gbuff[9][6] ,
         \gbuff[9][5] , \gbuff[9][4] , \gbuff[9][3] , \gbuff[9][2] ,
         \gbuff[9][1] , \gbuff[9][0] , \gbuff[8][31] , \gbuff[8][30] ,
         \gbuff[8][29] , \gbuff[8][28] , \gbuff[8][27] , \gbuff[8][26] ,
         \gbuff[8][25] , \gbuff[8][24] , \gbuff[8][23] , \gbuff[8][22] ,
         \gbuff[8][21] , \gbuff[8][20] , \gbuff[8][19] , \gbuff[8][18] ,
         \gbuff[8][17] , \gbuff[8][16] , \gbuff[8][15] , \gbuff[8][14] ,
         \gbuff[8][13] , \gbuff[8][12] , \gbuff[8][11] , \gbuff[8][10] ,
         \gbuff[8][9] , \gbuff[8][8] , \gbuff[8][7] , \gbuff[8][6] ,
         \gbuff[8][5] , \gbuff[8][4] , \gbuff[8][3] , \gbuff[8][2] ,
         \gbuff[8][1] , \gbuff[8][0] , \gbuff[11][31] , \gbuff[11][30] ,
         \gbuff[11][29] , \gbuff[11][28] , \gbuff[11][27] , \gbuff[11][26] ,
         \gbuff[11][25] , \gbuff[11][24] , \gbuff[11][23] , \gbuff[11][22] ,
         \gbuff[11][21] , \gbuff[11][20] , \gbuff[11][19] , \gbuff[11][18] ,
         \gbuff[11][17] , \gbuff[11][16] , \gbuff[11][15] , \gbuff[11][14] ,
         \gbuff[11][13] , \gbuff[11][12] , \gbuff[11][11] , \gbuff[11][10] ,
         \gbuff[11][9] , \gbuff[11][8] , \gbuff[11][7] , \gbuff[11][6] ,
         \gbuff[11][5] , \gbuff[11][4] , \gbuff[11][3] , \gbuff[11][2] ,
         \gbuff[11][1] , \gbuff[11][0] , \gbuff[10][31] , \gbuff[10][30] ,
         \gbuff[10][29] , \gbuff[10][28] , \gbuff[10][27] , \gbuff[10][26] ,
         \gbuff[10][25] , \gbuff[10][24] , \gbuff[10][23] , \gbuff[10][22] ,
         \gbuff[10][21] , \gbuff[10][20] , \gbuff[10][19] , \gbuff[10][18] ,
         \gbuff[10][17] , \gbuff[10][16] , \gbuff[10][15] , \gbuff[10][14] ,
         \gbuff[10][13] , \gbuff[10][12] , \gbuff[10][11] , \gbuff[10][10] ,
         \gbuff[10][9] , \gbuff[10][8] , \gbuff[10][7] , \gbuff[10][6] ,
         \gbuff[10][5] , \gbuff[10][4] , \gbuff[10][3] , \gbuff[10][2] ,
         \gbuff[10][1] , \gbuff[10][0] , \gbuff[13][31] , \gbuff[13][30] ,
         \gbuff[13][29] , \gbuff[13][28] , \gbuff[13][27] , \gbuff[13][26] ,
         \gbuff[13][25] , \gbuff[13][24] , \gbuff[13][23] , \gbuff[13][22] ,
         \gbuff[13][21] , \gbuff[13][20] , \gbuff[13][19] , \gbuff[13][18] ,
         \gbuff[13][17] , \gbuff[13][16] , \gbuff[13][15] , \gbuff[13][14] ,
         \gbuff[13][13] , \gbuff[13][12] , \gbuff[13][11] , \gbuff[13][10] ,
         \gbuff[13][9] , \gbuff[13][8] , \gbuff[13][7] , \gbuff[13][6] ,
         \gbuff[13][5] , \gbuff[13][4] , \gbuff[13][3] , \gbuff[13][2] ,
         \gbuff[13][1] , \gbuff[13][0] , \gbuff[12][31] , \gbuff[12][30] ,
         \gbuff[12][29] , \gbuff[12][28] , \gbuff[12][27] , \gbuff[12][26] ,
         \gbuff[12][25] , \gbuff[12][24] , \gbuff[12][23] , \gbuff[12][22] ,
         \gbuff[12][21] , \gbuff[12][20] , \gbuff[12][19] , \gbuff[12][18] ,
         \gbuff[12][17] , \gbuff[12][16] , \gbuff[12][15] , \gbuff[12][14] ,
         \gbuff[12][13] , \gbuff[12][12] , \gbuff[12][11] , \gbuff[12][10] ,
         \gbuff[12][9] , \gbuff[12][8] , \gbuff[12][7] , \gbuff[12][6] ,
         \gbuff[12][5] , \gbuff[12][4] , \gbuff[12][3] , \gbuff[12][2] ,
         \gbuff[12][1] , \gbuff[12][0] , \gbuff[15][31] , \gbuff[15][30] ,
         \gbuff[15][29] , \gbuff[15][28] , \gbuff[15][27] , \gbuff[15][26] ,
         \gbuff[15][25] , \gbuff[15][24] , \gbuff[15][23] , \gbuff[15][22] ,
         \gbuff[15][21] , \gbuff[15][20] , \gbuff[15][19] , \gbuff[15][18] ,
         \gbuff[15][17] , \gbuff[15][16] , \gbuff[15][15] , \gbuff[15][14] ,
         \gbuff[15][13] , \gbuff[15][12] , \gbuff[15][11] , \gbuff[15][10] ,
         \gbuff[15][9] , \gbuff[15][8] , \gbuff[15][7] , \gbuff[15][6] ,
         \gbuff[15][5] , \gbuff[15][4] , \gbuff[15][3] , \gbuff[15][2] ,
         \gbuff[15][1] , \gbuff[15][0] , \gbuff[14][31] , \gbuff[14][30] ,
         \gbuff[14][29] , \gbuff[14][28] , \gbuff[14][27] , \gbuff[14][26] ,
         \gbuff[14][25] , \gbuff[14][24] , \gbuff[14][23] , \gbuff[14][22] ,
         \gbuff[14][21] , \gbuff[14][20] , \gbuff[14][19] , \gbuff[14][18] ,
         \gbuff[14][17] , \gbuff[14][16] , \gbuff[14][15] , \gbuff[14][14] ,
         \gbuff[14][13] , \gbuff[14][12] , \gbuff[14][11] , \gbuff[14][10] ,
         \gbuff[14][9] , \gbuff[14][8] , \gbuff[14][7] , \gbuff[14][6] ,
         \gbuff[14][5] , \gbuff[14][4] , \gbuff[14][3] , \gbuff[14][2] ,
         \gbuff[14][1] , \gbuff[14][0] , \gbuff[17][31] , \gbuff[17][30] ,
         \gbuff[17][29] , \gbuff[17][28] , \gbuff[17][27] , \gbuff[17][26] ,
         \gbuff[17][25] , \gbuff[17][24] , \gbuff[17][23] , \gbuff[17][22] ,
         \gbuff[17][21] , \gbuff[17][20] , \gbuff[17][19] , \gbuff[17][18] ,
         \gbuff[17][17] , \gbuff[17][16] , \gbuff[17][15] , \gbuff[17][14] ,
         \gbuff[17][13] , \gbuff[17][12] , \gbuff[17][11] , \gbuff[17][10] ,
         \gbuff[17][9] , \gbuff[17][8] , \gbuff[17][7] , \gbuff[17][6] ,
         \gbuff[17][5] , \gbuff[17][4] , \gbuff[17][3] , \gbuff[17][2] ,
         \gbuff[17][1] , \gbuff[17][0] , \gbuff[16][31] , \gbuff[16][30] ,
         \gbuff[16][29] , \gbuff[16][28] , \gbuff[16][27] , \gbuff[16][26] ,
         \gbuff[16][25] , \gbuff[16][24] , \gbuff[16][23] , \gbuff[16][22] ,
         \gbuff[16][21] , \gbuff[16][20] , \gbuff[16][19] , \gbuff[16][18] ,
         \gbuff[16][17] , \gbuff[16][16] , \gbuff[16][15] , \gbuff[16][14] ,
         \gbuff[16][13] , \gbuff[16][12] , \gbuff[16][11] , \gbuff[16][10] ,
         \gbuff[16][9] , \gbuff[16][8] , \gbuff[16][7] , \gbuff[16][6] ,
         \gbuff[16][5] , \gbuff[16][4] , \gbuff[16][3] , \gbuff[16][2] ,
         \gbuff[16][1] , \gbuff[16][0] , \gbuff[19][31] , \gbuff[19][30] ,
         \gbuff[19][29] , \gbuff[19][28] , \gbuff[19][27] , \gbuff[19][26] ,
         \gbuff[19][25] , \gbuff[19][24] , \gbuff[19][23] , \gbuff[19][22] ,
         \gbuff[19][21] , \gbuff[19][20] , \gbuff[19][19] , \gbuff[19][18] ,
         \gbuff[19][17] , \gbuff[19][16] , \gbuff[19][15] , \gbuff[19][14] ,
         \gbuff[19][13] , \gbuff[19][12] , \gbuff[19][11] , \gbuff[19][10] ,
         \gbuff[19][9] , \gbuff[19][8] , \gbuff[19][7] , \gbuff[19][6] ,
         \gbuff[19][5] , \gbuff[19][4] , \gbuff[19][3] , \gbuff[19][2] ,
         \gbuff[19][1] , \gbuff[19][0] , \gbuff[18][31] , \gbuff[18][30] ,
         \gbuff[18][29] , \gbuff[18][28] , \gbuff[18][27] , \gbuff[18][26] ,
         \gbuff[18][25] , \gbuff[18][24] , \gbuff[18][23] , \gbuff[18][22] ,
         \gbuff[18][21] , \gbuff[18][20] , \gbuff[18][19] , \gbuff[18][18] ,
         \gbuff[18][17] , \gbuff[18][16] , \gbuff[18][15] , \gbuff[18][14] ,
         \gbuff[18][13] , \gbuff[18][12] , \gbuff[18][11] , \gbuff[18][10] ,
         \gbuff[18][9] , \gbuff[18][8] , \gbuff[18][7] , \gbuff[18][6] ,
         \gbuff[18][5] , \gbuff[18][4] , \gbuff[18][3] , \gbuff[18][2] ,
         \gbuff[18][1] , \gbuff[18][0] , \gbuff[21][31] , \gbuff[21][30] ,
         \gbuff[21][29] , \gbuff[21][28] , \gbuff[21][27] , \gbuff[21][26] ,
         \gbuff[21][25] , \gbuff[21][24] , \gbuff[21][23] , \gbuff[21][22] ,
         \gbuff[21][21] , \gbuff[21][20] , \gbuff[21][19] , \gbuff[21][18] ,
         \gbuff[21][17] , \gbuff[21][16] , \gbuff[21][15] , \gbuff[21][14] ,
         \gbuff[21][13] , \gbuff[21][12] , \gbuff[21][11] , \gbuff[21][10] ,
         \gbuff[21][9] , \gbuff[21][8] , \gbuff[21][7] , \gbuff[21][6] ,
         \gbuff[21][5] , \gbuff[21][4] , \gbuff[21][3] , \gbuff[21][2] ,
         \gbuff[21][1] , \gbuff[21][0] , \gbuff[20][31] , \gbuff[20][30] ,
         \gbuff[20][29] , \gbuff[20][28] , \gbuff[20][27] , \gbuff[20][26] ,
         \gbuff[20][25] , \gbuff[20][24] , \gbuff[20][23] , \gbuff[20][22] ,
         \gbuff[20][21] , \gbuff[20][20] , \gbuff[20][19] , \gbuff[20][18] ,
         \gbuff[20][17] , \gbuff[20][16] , \gbuff[20][15] , \gbuff[20][14] ,
         \gbuff[20][13] , \gbuff[20][12] , \gbuff[20][11] , \gbuff[20][10] ,
         \gbuff[20][9] , \gbuff[20][8] , \gbuff[20][7] , \gbuff[20][6] ,
         \gbuff[20][5] , \gbuff[20][4] , \gbuff[20][3] , \gbuff[20][2] ,
         \gbuff[20][1] , \gbuff[20][0] , \gbuff[23][31] , \gbuff[23][30] ,
         \gbuff[23][29] , \gbuff[23][28] , \gbuff[23][27] , \gbuff[23][26] ,
         \gbuff[23][25] , \gbuff[23][24] , \gbuff[23][23] , \gbuff[23][22] ,
         \gbuff[23][21] , \gbuff[23][20] , \gbuff[23][19] , \gbuff[23][18] ,
         \gbuff[23][17] , \gbuff[23][16] , \gbuff[23][15] , \gbuff[23][14] ,
         \gbuff[23][13] , \gbuff[23][12] , \gbuff[23][11] , \gbuff[23][10] ,
         \gbuff[23][9] , \gbuff[23][8] , \gbuff[23][7] , \gbuff[23][6] ,
         \gbuff[23][5] , \gbuff[23][4] , \gbuff[23][3] , \gbuff[23][2] ,
         \gbuff[23][1] , \gbuff[23][0] , \gbuff[22][31] , \gbuff[22][30] ,
         \gbuff[22][29] , \gbuff[22][28] , \gbuff[22][27] , \gbuff[22][26] ,
         \gbuff[22][25] , \gbuff[22][24] , \gbuff[22][23] , \gbuff[22][22] ,
         \gbuff[22][21] , \gbuff[22][20] , \gbuff[22][19] , \gbuff[22][18] ,
         \gbuff[22][17] , \gbuff[22][16] , \gbuff[22][15] , \gbuff[22][14] ,
         \gbuff[22][13] , \gbuff[22][12] , \gbuff[22][11] , \gbuff[22][10] ,
         \gbuff[22][9] , \gbuff[22][8] , \gbuff[22][7] , \gbuff[22][6] ,
         \gbuff[22][5] , \gbuff[22][4] , \gbuff[22][3] , \gbuff[22][2] ,
         \gbuff[22][1] , \gbuff[22][0] , \gbuff[25][31] , \gbuff[25][30] ,
         \gbuff[25][29] , \gbuff[25][28] , \gbuff[25][27] , \gbuff[25][26] ,
         \gbuff[25][25] , \gbuff[25][24] , \gbuff[25][23] , \gbuff[25][22] ,
         \gbuff[25][21] , \gbuff[25][20] , \gbuff[25][19] , \gbuff[25][18] ,
         \gbuff[25][17] , \gbuff[25][16] , \gbuff[25][15] , \gbuff[25][14] ,
         \gbuff[25][13] , \gbuff[25][12] , \gbuff[25][11] , \gbuff[25][10] ,
         \gbuff[25][9] , \gbuff[25][8] , \gbuff[25][7] , \gbuff[25][6] ,
         \gbuff[25][5] , \gbuff[25][4] , \gbuff[25][3] , \gbuff[25][2] ,
         \gbuff[25][1] , \gbuff[25][0] , \gbuff[24][31] , \gbuff[24][30] ,
         \gbuff[24][29] , \gbuff[24][28] , \gbuff[24][27] , \gbuff[24][26] ,
         \gbuff[24][25] , \gbuff[24][24] , \gbuff[24][23] , \gbuff[24][22] ,
         \gbuff[24][21] , \gbuff[24][20] , \gbuff[24][19] , \gbuff[24][18] ,
         \gbuff[24][17] , \gbuff[24][16] , \gbuff[24][15] , \gbuff[24][14] ,
         \gbuff[24][13] , \gbuff[24][12] , \gbuff[24][11] , \gbuff[24][10] ,
         \gbuff[24][9] , \gbuff[24][8] , \gbuff[24][7] , \gbuff[24][6] ,
         \gbuff[24][5] , \gbuff[24][4] , \gbuff[24][3] , \gbuff[24][2] ,
         \gbuff[24][1] , \gbuff[24][0] , \gbuff[27][31] , \gbuff[27][30] ,
         \gbuff[27][29] , \gbuff[27][28] , \gbuff[27][27] , \gbuff[27][26] ,
         \gbuff[27][25] , \gbuff[27][24] , \gbuff[27][23] , \gbuff[27][22] ,
         \gbuff[27][21] , \gbuff[27][20] , \gbuff[27][19] , \gbuff[27][18] ,
         \gbuff[27][17] , \gbuff[27][16] , \gbuff[27][15] , \gbuff[27][14] ,
         \gbuff[27][13] , \gbuff[27][12] , \gbuff[27][11] , \gbuff[27][10] ,
         \gbuff[27][9] , \gbuff[27][8] , \gbuff[27][7] , \gbuff[27][6] ,
         \gbuff[27][5] , \gbuff[27][4] , \gbuff[27][3] , \gbuff[27][2] ,
         \gbuff[27][1] , \gbuff[27][0] , \gbuff[26][31] , \gbuff[26][30] ,
         \gbuff[26][29] , \gbuff[26][28] , \gbuff[26][27] , \gbuff[26][26] ,
         \gbuff[26][25] , \gbuff[26][24] , \gbuff[26][23] , \gbuff[26][22] ,
         \gbuff[26][21] , \gbuff[26][20] , \gbuff[26][19] , \gbuff[26][18] ,
         \gbuff[26][17] , \gbuff[26][16] , \gbuff[26][15] , \gbuff[26][14] ,
         \gbuff[26][13] , \gbuff[26][12] , \gbuff[26][11] , \gbuff[26][10] ,
         \gbuff[26][9] , \gbuff[26][8] , \gbuff[26][7] , \gbuff[26][6] ,
         \gbuff[26][5] , \gbuff[26][4] , \gbuff[26][3] , \gbuff[26][2] ,
         \gbuff[26][1] , \gbuff[26][0] , \gbuff[29][31] , \gbuff[29][30] ,
         \gbuff[29][29] , \gbuff[29][28] , \gbuff[29][27] , \gbuff[29][26] ,
         \gbuff[29][25] , \gbuff[29][24] , \gbuff[29][23] , \gbuff[29][22] ,
         \gbuff[29][21] , \gbuff[29][20] , \gbuff[29][19] , \gbuff[29][18] ,
         \gbuff[29][17] , \gbuff[29][16] , \gbuff[29][15] , \gbuff[29][14] ,
         \gbuff[29][13] , \gbuff[29][12] , \gbuff[29][11] , \gbuff[29][10] ,
         \gbuff[29][9] , \gbuff[29][8] , \gbuff[29][7] , \gbuff[29][6] ,
         \gbuff[29][5] , \gbuff[29][4] , \gbuff[29][3] , \gbuff[29][2] ,
         \gbuff[29][1] , \gbuff[29][0] , \gbuff[28][31] , \gbuff[28][30] ,
         \gbuff[28][29] , \gbuff[28][28] , \gbuff[28][27] , \gbuff[28][26] ,
         \gbuff[28][25] , \gbuff[28][24] , \gbuff[28][23] , \gbuff[28][22] ,
         \gbuff[28][21] , \gbuff[28][20] , \gbuff[28][19] , \gbuff[28][18] ,
         \gbuff[28][17] , \gbuff[28][16] , \gbuff[28][15] , \gbuff[28][14] ,
         \gbuff[28][13] , \gbuff[28][12] , \gbuff[28][11] , \gbuff[28][10] ,
         \gbuff[28][9] , \gbuff[28][8] , \gbuff[28][7] , \gbuff[28][6] ,
         \gbuff[28][5] , \gbuff[28][4] , \gbuff[28][3] , \gbuff[28][2] ,
         \gbuff[28][1] , \gbuff[28][0] , \gbuff[31][31] , \gbuff[31][30] ,
         \gbuff[31][29] , \gbuff[31][28] , \gbuff[31][27] , \gbuff[31][26] ,
         \gbuff[31][25] , \gbuff[31][24] , \gbuff[31][23] , \gbuff[31][22] ,
         \gbuff[31][21] , \gbuff[31][20] , \gbuff[31][19] , \gbuff[31][18] ,
         \gbuff[31][17] , \gbuff[31][16] , \gbuff[31][15] , \gbuff[31][14] ,
         \gbuff[31][13] , \gbuff[31][12] , \gbuff[31][11] , \gbuff[31][10] ,
         \gbuff[31][9] , \gbuff[31][8] , \gbuff[31][7] , \gbuff[31][6] ,
         \gbuff[31][5] , \gbuff[31][4] , \gbuff[31][3] , \gbuff[31][2] ,
         \gbuff[31][1] , \gbuff[31][0] , \gbuff[30][31] , \gbuff[30][30] ,
         \gbuff[30][29] , \gbuff[30][28] , \gbuff[30][27] , \gbuff[30][26] ,
         \gbuff[30][25] , \gbuff[30][24] , \gbuff[30][23] , \gbuff[30][22] ,
         \gbuff[30][21] , \gbuff[30][20] , \gbuff[30][19] , \gbuff[30][18] ,
         \gbuff[30][17] , \gbuff[30][16] , \gbuff[30][15] , \gbuff[30][14] ,
         \gbuff[30][13] , \gbuff[30][12] , \gbuff[30][11] , \gbuff[30][10] ,
         \gbuff[30][9] , \gbuff[30][8] , \gbuff[30][7] , \gbuff[30][6] ,
         \gbuff[30][5] , \gbuff[30][4] , \gbuff[30][3] , \gbuff[30][2] ,
         \gbuff[30][1] , \gbuff[30][0] , N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N81, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n104, n106, n108, n110, n112, n114, n116, n119, n121, n122,
         n123, n124, n125, n126, n127, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824;
  assign N10 = index[0];
  assign N11 = index[1];
  assign N12 = index[2];
  assign N13 = index[3];
  assign N14 = index[4];

  DFFRX1 \gbuff_reg[29][31]  ( .D(n1836), .CK(clk), .RN(n1521), .Q(
        \gbuff[29][31] ) );
  DFFRX1 \gbuff_reg[29][30]  ( .D(n1837), .CK(clk), .RN(n1521), .Q(
        \gbuff[29][30] ) );
  DFFRX1 \gbuff_reg[29][29]  ( .D(n1838), .CK(clk), .RN(n1521), .Q(
        \gbuff[29][29] ) );
  DFFRX1 \gbuff_reg[29][28]  ( .D(n1839), .CK(clk), .RN(n1521), .Q(
        \gbuff[29][28] ) );
  DFFRX1 \gbuff_reg[29][27]  ( .D(n1840), .CK(clk), .RN(n1521), .Q(
        \gbuff[29][27] ) );
  DFFRX1 \gbuff_reg[29][26]  ( .D(n1841), .CK(clk), .RN(n1521), .Q(
        \gbuff[29][26] ) );
  DFFRX1 \gbuff_reg[29][25]  ( .D(n1842), .CK(clk), .RN(n1521), .Q(
        \gbuff[29][25] ) );
  DFFRX1 \gbuff_reg[29][24]  ( .D(n1843), .CK(clk), .RN(n1521), .Q(
        \gbuff[29][24] ) );
  DFFRX1 \gbuff_reg[29][23]  ( .D(n1844), .CK(clk), .RN(n1521), .Q(
        \gbuff[29][23] ) );
  DFFRX1 \gbuff_reg[29][22]  ( .D(n1845), .CK(clk), .RN(n1521), .Q(
        \gbuff[29][22] ) );
  DFFRX1 \gbuff_reg[29][21]  ( .D(n1846), .CK(clk), .RN(n1521), .Q(
        \gbuff[29][21] ) );
  DFFRX1 \gbuff_reg[29][20]  ( .D(n1847), .CK(clk), .RN(n1521), .Q(
        \gbuff[29][20] ) );
  DFFRX1 \gbuff_reg[29][19]  ( .D(n1848), .CK(clk), .RN(n1520), .Q(
        \gbuff[29][19] ) );
  DFFRX1 \gbuff_reg[29][18]  ( .D(n1849), .CK(clk), .RN(n1520), .Q(
        \gbuff[29][18] ) );
  DFFRX1 \gbuff_reg[29][17]  ( .D(n1850), .CK(clk), .RN(n1520), .Q(
        \gbuff[29][17] ) );
  DFFRX1 \gbuff_reg[29][16]  ( .D(n1851), .CK(clk), .RN(n1520), .Q(
        \gbuff[29][16] ) );
  DFFRX1 \gbuff_reg[29][15]  ( .D(n1852), .CK(clk), .RN(n1520), .Q(
        \gbuff[29][15] ) );
  DFFRX1 \gbuff_reg[29][14]  ( .D(n1853), .CK(clk), .RN(n1520), .Q(
        \gbuff[29][14] ) );
  DFFRX1 \gbuff_reg[29][13]  ( .D(n1854), .CK(clk), .RN(n1520), .Q(
        \gbuff[29][13] ) );
  DFFRX1 \gbuff_reg[29][12]  ( .D(n1855), .CK(clk), .RN(n1520), .Q(
        \gbuff[29][12] ) );
  DFFRX1 \gbuff_reg[29][11]  ( .D(n1856), .CK(clk), .RN(n1520), .Q(
        \gbuff[29][11] ) );
  DFFRX1 \gbuff_reg[29][10]  ( .D(n1857), .CK(clk), .RN(n1520), .Q(
        \gbuff[29][10] ) );
  DFFRX1 \gbuff_reg[29][9]  ( .D(n1858), .CK(clk), .RN(n1520), .Q(
        \gbuff[29][9] ) );
  DFFRX1 \gbuff_reg[29][8]  ( .D(n1859), .CK(clk), .RN(n1520), .Q(
        \gbuff[29][8] ) );
  DFFRX1 \gbuff_reg[29][7]  ( .D(n1860), .CK(clk), .RN(n1519), .Q(
        \gbuff[29][7] ) );
  DFFRX1 \gbuff_reg[29][6]  ( .D(n1861), .CK(clk), .RN(n1519), .Q(
        \gbuff[29][6] ) );
  DFFRX1 \gbuff_reg[29][5]  ( .D(n1862), .CK(clk), .RN(n1519), .Q(
        \gbuff[29][5] ) );
  DFFRX1 \gbuff_reg[29][4]  ( .D(n1863), .CK(clk), .RN(n1519), .Q(
        \gbuff[29][4] ) );
  DFFRX1 \gbuff_reg[29][3]  ( .D(n1864), .CK(clk), .RN(n1519), .Q(
        \gbuff[29][3] ) );
  DFFRX1 \gbuff_reg[29][2]  ( .D(n1865), .CK(clk), .RN(n1519), .Q(
        \gbuff[29][2] ) );
  DFFRX1 \gbuff_reg[29][1]  ( .D(n1866), .CK(clk), .RN(n1519), .Q(
        \gbuff[29][1] ) );
  DFFRX1 \gbuff_reg[29][0]  ( .D(n1867), .CK(clk), .RN(n1519), .Q(
        \gbuff[29][0] ) );
  DFFRX1 \gbuff_reg[25][31]  ( .D(n1964), .CK(clk), .RN(n1511), .Q(
        \gbuff[25][31] ) );
  DFFRX1 \gbuff_reg[25][30]  ( .D(n1965), .CK(clk), .RN(n1511), .Q(
        \gbuff[25][30] ) );
  DFFRX1 \gbuff_reg[25][29]  ( .D(n1966), .CK(clk), .RN(n1511), .Q(
        \gbuff[25][29] ) );
  DFFRX1 \gbuff_reg[25][28]  ( .D(n1967), .CK(clk), .RN(n1511), .Q(
        \gbuff[25][28] ) );
  DFFRX1 \gbuff_reg[25][27]  ( .D(n1968), .CK(clk), .RN(n1510), .Q(
        \gbuff[25][27] ) );
  DFFRX1 \gbuff_reg[25][26]  ( .D(n1969), .CK(clk), .RN(n1510), .Q(
        \gbuff[25][26] ) );
  DFFRX1 \gbuff_reg[25][25]  ( .D(n1970), .CK(clk), .RN(n1510), .Q(
        \gbuff[25][25] ) );
  DFFRX1 \gbuff_reg[25][24]  ( .D(n1971), .CK(clk), .RN(n1510), .Q(
        \gbuff[25][24] ) );
  DFFRX1 \gbuff_reg[25][23]  ( .D(n1972), .CK(clk), .RN(n1510), .Q(
        \gbuff[25][23] ) );
  DFFRX1 \gbuff_reg[25][22]  ( .D(n1973), .CK(clk), .RN(n1510), .Q(
        \gbuff[25][22] ) );
  DFFRX1 \gbuff_reg[25][21]  ( .D(n1974), .CK(clk), .RN(n1510), .Q(
        \gbuff[25][21] ) );
  DFFRX1 \gbuff_reg[25][20]  ( .D(n1975), .CK(clk), .RN(n1510), .Q(
        \gbuff[25][20] ) );
  DFFRX1 \gbuff_reg[25][19]  ( .D(n1976), .CK(clk), .RN(n1510), .Q(
        \gbuff[25][19] ) );
  DFFRX1 \gbuff_reg[25][18]  ( .D(n1977), .CK(clk), .RN(n1510), .Q(
        \gbuff[25][18] ) );
  DFFRX1 \gbuff_reg[25][17]  ( .D(n1978), .CK(clk), .RN(n1510), .Q(
        \gbuff[25][17] ) );
  DFFRX1 \gbuff_reg[25][16]  ( .D(n1979), .CK(clk), .RN(n1510), .Q(
        \gbuff[25][16] ) );
  DFFRX1 \gbuff_reg[25][15]  ( .D(n1980), .CK(clk), .RN(n1509), .Q(
        \gbuff[25][15] ) );
  DFFRX1 \gbuff_reg[25][14]  ( .D(n1981), .CK(clk), .RN(n1509), .Q(
        \gbuff[25][14] ) );
  DFFRX1 \gbuff_reg[25][13]  ( .D(n1982), .CK(clk), .RN(n1509), .Q(
        \gbuff[25][13] ) );
  DFFRX1 \gbuff_reg[25][12]  ( .D(n1983), .CK(clk), .RN(n1509), .Q(
        \gbuff[25][12] ) );
  DFFRX1 \gbuff_reg[25][11]  ( .D(n1984), .CK(clk), .RN(n1509), .Q(
        \gbuff[25][11] ) );
  DFFRX1 \gbuff_reg[25][10]  ( .D(n1985), .CK(clk), .RN(n1509), .Q(
        \gbuff[25][10] ) );
  DFFRX1 \gbuff_reg[25][9]  ( .D(n1986), .CK(clk), .RN(n1509), .Q(
        \gbuff[25][9] ) );
  DFFRX1 \gbuff_reg[25][8]  ( .D(n1987), .CK(clk), .RN(n1509), .Q(
        \gbuff[25][8] ) );
  DFFRX1 \gbuff_reg[25][7]  ( .D(n1988), .CK(clk), .RN(n1509), .Q(
        \gbuff[25][7] ) );
  DFFRX1 \gbuff_reg[25][6]  ( .D(n1989), .CK(clk), .RN(n1509), .Q(
        \gbuff[25][6] ) );
  DFFRX1 \gbuff_reg[25][5]  ( .D(n1990), .CK(clk), .RN(n1509), .Q(
        \gbuff[25][5] ) );
  DFFRX1 \gbuff_reg[25][4]  ( .D(n1991), .CK(clk), .RN(n1509), .Q(
        \gbuff[25][4] ) );
  DFFRX1 \gbuff_reg[25][3]  ( .D(n1992), .CK(clk), .RN(n1508), .Q(
        \gbuff[25][3] ) );
  DFFRX1 \gbuff_reg[25][2]  ( .D(n1993), .CK(clk), .RN(n1508), .Q(
        \gbuff[25][2] ) );
  DFFRX1 \gbuff_reg[25][1]  ( .D(n1994), .CK(clk), .RN(n1508), .Q(
        \gbuff[25][1] ) );
  DFFRX1 \gbuff_reg[25][0]  ( .D(n1995), .CK(clk), .RN(n1508), .Q(
        \gbuff[25][0] ) );
  DFFRX1 \gbuff_reg[21][31]  ( .D(n2092), .CK(clk), .RN(n1500), .Q(
        \gbuff[21][31] ) );
  DFFRX1 \gbuff_reg[21][30]  ( .D(n2093), .CK(clk), .RN(n1500), .Q(
        \gbuff[21][30] ) );
  DFFRX1 \gbuff_reg[21][29]  ( .D(n2094), .CK(clk), .RN(n1500), .Q(
        \gbuff[21][29] ) );
  DFFRX1 \gbuff_reg[21][28]  ( .D(n2095), .CK(clk), .RN(n1500), .Q(
        \gbuff[21][28] ) );
  DFFRX1 \gbuff_reg[21][27]  ( .D(n2096), .CK(clk), .RN(n1500), .Q(
        \gbuff[21][27] ) );
  DFFRX1 \gbuff_reg[21][26]  ( .D(n2097), .CK(clk), .RN(n1500), .Q(
        \gbuff[21][26] ) );
  DFFRX1 \gbuff_reg[21][25]  ( .D(n2098), .CK(clk), .RN(n1500), .Q(
        \gbuff[21][25] ) );
  DFFRX1 \gbuff_reg[21][24]  ( .D(n2099), .CK(clk), .RN(n1500), .Q(
        \gbuff[21][24] ) );
  DFFRX1 \gbuff_reg[21][23]  ( .D(n2100), .CK(clk), .RN(n1499), .Q(
        \gbuff[21][23] ) );
  DFFRX1 \gbuff_reg[21][22]  ( .D(n2101), .CK(clk), .RN(n1499), .Q(
        \gbuff[21][22] ) );
  DFFRX1 \gbuff_reg[21][21]  ( .D(n2102), .CK(clk), .RN(n1499), .Q(
        \gbuff[21][21] ) );
  DFFRX1 \gbuff_reg[21][20]  ( .D(n2103), .CK(clk), .RN(n1499), .Q(
        \gbuff[21][20] ) );
  DFFRX1 \gbuff_reg[21][19]  ( .D(n2104), .CK(clk), .RN(n1499), .Q(
        \gbuff[21][19] ) );
  DFFRX1 \gbuff_reg[21][18]  ( .D(n2105), .CK(clk), .RN(n1499), .Q(
        \gbuff[21][18] ) );
  DFFRX1 \gbuff_reg[21][17]  ( .D(n2106), .CK(clk), .RN(n1499), .Q(
        \gbuff[21][17] ) );
  DFFRX1 \gbuff_reg[21][16]  ( .D(n2107), .CK(clk), .RN(n1499), .Q(
        \gbuff[21][16] ) );
  DFFRX1 \gbuff_reg[21][15]  ( .D(n2108), .CK(clk), .RN(n1499), .Q(
        \gbuff[21][15] ) );
  DFFRX1 \gbuff_reg[21][14]  ( .D(n2109), .CK(clk), .RN(n1499), .Q(
        \gbuff[21][14] ) );
  DFFRX1 \gbuff_reg[21][13]  ( .D(n2110), .CK(clk), .RN(n1499), .Q(
        \gbuff[21][13] ) );
  DFFRX1 \gbuff_reg[21][12]  ( .D(n2111), .CK(clk), .RN(n1499), .Q(
        \gbuff[21][12] ) );
  DFFRX1 \gbuff_reg[21][11]  ( .D(n2112), .CK(clk), .RN(n1498), .Q(
        \gbuff[21][11] ) );
  DFFRX1 \gbuff_reg[21][10]  ( .D(n2113), .CK(clk), .RN(n1498), .Q(
        \gbuff[21][10] ) );
  DFFRX1 \gbuff_reg[21][9]  ( .D(n2114), .CK(clk), .RN(n1498), .Q(
        \gbuff[21][9] ) );
  DFFRX1 \gbuff_reg[21][8]  ( .D(n2115), .CK(clk), .RN(n1498), .Q(
        \gbuff[21][8] ) );
  DFFRX1 \gbuff_reg[21][7]  ( .D(n2116), .CK(clk), .RN(n1498), .Q(
        \gbuff[21][7] ) );
  DFFRX1 \gbuff_reg[21][6]  ( .D(n2117), .CK(clk), .RN(n1498), .Q(
        \gbuff[21][6] ) );
  DFFRX1 \gbuff_reg[21][5]  ( .D(n2118), .CK(clk), .RN(n1498), .Q(
        \gbuff[21][5] ) );
  DFFRX1 \gbuff_reg[21][4]  ( .D(n2119), .CK(clk), .RN(n1498), .Q(
        \gbuff[21][4] ) );
  DFFRX1 \gbuff_reg[21][3]  ( .D(n2120), .CK(clk), .RN(n1498), .Q(
        \gbuff[21][3] ) );
  DFFRX1 \gbuff_reg[21][2]  ( .D(n2121), .CK(clk), .RN(n1498), .Q(
        \gbuff[21][2] ) );
  DFFRX1 \gbuff_reg[21][1]  ( .D(n2122), .CK(clk), .RN(n1498), .Q(
        \gbuff[21][1] ) );
  DFFRX1 \gbuff_reg[21][0]  ( .D(n2123), .CK(clk), .RN(n1498), .Q(
        \gbuff[21][0] ) );
  DFFRX1 \gbuff_reg[17][31]  ( .D(n2220), .CK(clk), .RN(n1489), .Q(
        \gbuff[17][31] ) );
  DFFRX1 \gbuff_reg[17][30]  ( .D(n2221), .CK(clk), .RN(n1489), .Q(
        \gbuff[17][30] ) );
  DFFRX1 \gbuff_reg[17][29]  ( .D(n2222), .CK(clk), .RN(n1489), .Q(
        \gbuff[17][29] ) );
  DFFRX1 \gbuff_reg[17][28]  ( .D(n2223), .CK(clk), .RN(n1489), .Q(
        \gbuff[17][28] ) );
  DFFRX1 \gbuff_reg[17][27]  ( .D(n2224), .CK(clk), .RN(n1489), .Q(
        \gbuff[17][27] ) );
  DFFRX1 \gbuff_reg[17][26]  ( .D(n2225), .CK(clk), .RN(n1489), .Q(
        \gbuff[17][26] ) );
  DFFRX1 \gbuff_reg[17][25]  ( .D(n2226), .CK(clk), .RN(n1489), .Q(
        \gbuff[17][25] ) );
  DFFRX1 \gbuff_reg[17][24]  ( .D(n2227), .CK(clk), .RN(n1489), .Q(
        \gbuff[17][24] ) );
  DFFRX1 \gbuff_reg[17][23]  ( .D(n2228), .CK(clk), .RN(n1489), .Q(
        \gbuff[17][23] ) );
  DFFRX1 \gbuff_reg[17][22]  ( .D(n2229), .CK(clk), .RN(n1489), .Q(
        \gbuff[17][22] ) );
  DFFRX1 \gbuff_reg[17][21]  ( .D(n2230), .CK(clk), .RN(n1489), .Q(
        \gbuff[17][21] ) );
  DFFRX1 \gbuff_reg[17][20]  ( .D(n2231), .CK(clk), .RN(n1489), .Q(
        \gbuff[17][20] ) );
  DFFRX1 \gbuff_reg[17][19]  ( .D(n2232), .CK(clk), .RN(n1488), .Q(
        \gbuff[17][19] ) );
  DFFRX1 \gbuff_reg[17][18]  ( .D(n2233), .CK(clk), .RN(n1488), .Q(
        \gbuff[17][18] ) );
  DFFRX1 \gbuff_reg[17][17]  ( .D(n2234), .CK(clk), .RN(n1488), .Q(
        \gbuff[17][17] ) );
  DFFRX1 \gbuff_reg[17][16]  ( .D(n2235), .CK(clk), .RN(n1488), .Q(
        \gbuff[17][16] ) );
  DFFRX1 \gbuff_reg[17][15]  ( .D(n2236), .CK(clk), .RN(n1488), .Q(
        \gbuff[17][15] ) );
  DFFRX1 \gbuff_reg[17][14]  ( .D(n2237), .CK(clk), .RN(n1488), .Q(
        \gbuff[17][14] ) );
  DFFRX1 \gbuff_reg[17][13]  ( .D(n2238), .CK(clk), .RN(n1488), .Q(
        \gbuff[17][13] ) );
  DFFRX1 \gbuff_reg[17][12]  ( .D(n2239), .CK(clk), .RN(n1488), .Q(
        \gbuff[17][12] ) );
  DFFRX1 \gbuff_reg[17][11]  ( .D(n2240), .CK(clk), .RN(n1488), .Q(
        \gbuff[17][11] ) );
  DFFRX1 \gbuff_reg[17][10]  ( .D(n2241), .CK(clk), .RN(n1488), .Q(
        \gbuff[17][10] ) );
  DFFRX1 \gbuff_reg[17][9]  ( .D(n2242), .CK(clk), .RN(n1488), .Q(
        \gbuff[17][9] ) );
  DFFRX1 \gbuff_reg[17][8]  ( .D(n2243), .CK(clk), .RN(n1488), .Q(
        \gbuff[17][8] ) );
  DFFRX1 \gbuff_reg[17][7]  ( .D(n2244), .CK(clk), .RN(n1487), .Q(
        \gbuff[17][7] ) );
  DFFRX1 \gbuff_reg[17][6]  ( .D(n2245), .CK(clk), .RN(n1487), .Q(
        \gbuff[17][6] ) );
  DFFRX1 \gbuff_reg[17][5]  ( .D(n2246), .CK(clk), .RN(n1487), .Q(
        \gbuff[17][5] ) );
  DFFRX1 \gbuff_reg[17][4]  ( .D(n2247), .CK(clk), .RN(n1487), .Q(
        \gbuff[17][4] ) );
  DFFRX1 \gbuff_reg[17][3]  ( .D(n2248), .CK(clk), .RN(n1487), .Q(
        \gbuff[17][3] ) );
  DFFRX1 \gbuff_reg[17][2]  ( .D(n2249), .CK(clk), .RN(n1487), .Q(
        \gbuff[17][2] ) );
  DFFRX1 \gbuff_reg[17][1]  ( .D(n2250), .CK(clk), .RN(n1487), .Q(
        \gbuff[17][1] ) );
  DFFRX1 \gbuff_reg[17][0]  ( .D(n2251), .CK(clk), .RN(n1487), .Q(
        \gbuff[17][0] ) );
  DFFRX1 \gbuff_reg[13][31]  ( .D(n2348), .CK(clk), .RN(n1479), .Q(
        \gbuff[13][31] ) );
  DFFRX1 \gbuff_reg[13][30]  ( .D(n2349), .CK(clk), .RN(n1479), .Q(
        \gbuff[13][30] ) );
  DFFRX1 \gbuff_reg[13][29]  ( .D(n2350), .CK(clk), .RN(n1479), .Q(
        \gbuff[13][29] ) );
  DFFRX1 \gbuff_reg[13][28]  ( .D(n2351), .CK(clk), .RN(n1479), .Q(
        \gbuff[13][28] ) );
  DFFRX1 \gbuff_reg[13][27]  ( .D(n2352), .CK(clk), .RN(n1478), .Q(
        \gbuff[13][27] ) );
  DFFRX1 \gbuff_reg[13][26]  ( .D(n2353), .CK(clk), .RN(n1478), .Q(
        \gbuff[13][26] ) );
  DFFRX1 \gbuff_reg[13][25]  ( .D(n2354), .CK(clk), .RN(n1478), .Q(
        \gbuff[13][25] ) );
  DFFRX1 \gbuff_reg[13][24]  ( .D(n2355), .CK(clk), .RN(n1478), .Q(
        \gbuff[13][24] ) );
  DFFRX1 \gbuff_reg[13][23]  ( .D(n2356), .CK(clk), .RN(n1478), .Q(
        \gbuff[13][23] ) );
  DFFRX1 \gbuff_reg[13][22]  ( .D(n2357), .CK(clk), .RN(n1478), .Q(
        \gbuff[13][22] ) );
  DFFRX1 \gbuff_reg[13][21]  ( .D(n2358), .CK(clk), .RN(n1478), .Q(
        \gbuff[13][21] ) );
  DFFRX1 \gbuff_reg[13][20]  ( .D(n2359), .CK(clk), .RN(n1478), .Q(
        \gbuff[13][20] ) );
  DFFRX1 \gbuff_reg[13][19]  ( .D(n2360), .CK(clk), .RN(n1478), .Q(
        \gbuff[13][19] ) );
  DFFRX1 \gbuff_reg[13][18]  ( .D(n2361), .CK(clk), .RN(n1478), .Q(
        \gbuff[13][18] ) );
  DFFRX1 \gbuff_reg[13][17]  ( .D(n2362), .CK(clk), .RN(n1478), .Q(
        \gbuff[13][17] ) );
  DFFRX1 \gbuff_reg[13][16]  ( .D(n2363), .CK(clk), .RN(n1478), .Q(
        \gbuff[13][16] ) );
  DFFRX1 \gbuff_reg[13][15]  ( .D(n2364), .CK(clk), .RN(n1477), .Q(
        \gbuff[13][15] ) );
  DFFRX1 \gbuff_reg[13][14]  ( .D(n2365), .CK(clk), .RN(n1477), .Q(
        \gbuff[13][14] ) );
  DFFRX1 \gbuff_reg[13][13]  ( .D(n2366), .CK(clk), .RN(n1477), .Q(
        \gbuff[13][13] ) );
  DFFRX1 \gbuff_reg[13][12]  ( .D(n2367), .CK(clk), .RN(n1477), .Q(
        \gbuff[13][12] ) );
  DFFRX1 \gbuff_reg[13][11]  ( .D(n2368), .CK(clk), .RN(n1477), .Q(
        \gbuff[13][11] ) );
  DFFRX1 \gbuff_reg[13][10]  ( .D(n2369), .CK(clk), .RN(n1477), .Q(
        \gbuff[13][10] ) );
  DFFRX1 \gbuff_reg[13][9]  ( .D(n2370), .CK(clk), .RN(n1477), .Q(
        \gbuff[13][9] ) );
  DFFRX1 \gbuff_reg[13][8]  ( .D(n2371), .CK(clk), .RN(n1477), .Q(
        \gbuff[13][8] ) );
  DFFRX1 \gbuff_reg[13][7]  ( .D(n2372), .CK(clk), .RN(n1477), .Q(
        \gbuff[13][7] ) );
  DFFRX1 \gbuff_reg[13][6]  ( .D(n2373), .CK(clk), .RN(n1477), .Q(
        \gbuff[13][6] ) );
  DFFRX1 \gbuff_reg[13][5]  ( .D(n2374), .CK(clk), .RN(n1477), .Q(
        \gbuff[13][5] ) );
  DFFRX1 \gbuff_reg[13][4]  ( .D(n2375), .CK(clk), .RN(n1477), .Q(
        \gbuff[13][4] ) );
  DFFRX1 \gbuff_reg[13][3]  ( .D(n2376), .CK(clk), .RN(n1476), .Q(
        \gbuff[13][3] ) );
  DFFRX1 \gbuff_reg[13][2]  ( .D(n2377), .CK(clk), .RN(n1476), .Q(
        \gbuff[13][2] ) );
  DFFRX1 \gbuff_reg[13][1]  ( .D(n2378), .CK(clk), .RN(n1476), .Q(
        \gbuff[13][1] ) );
  DFFRX1 \gbuff_reg[13][0]  ( .D(n2379), .CK(clk), .RN(n1476), .Q(
        \gbuff[13][0] ) );
  DFFRX1 \gbuff_reg[9][31]  ( .D(n2476), .CK(clk), .RN(n1468), .Q(
        \gbuff[9][31] ) );
  DFFRX1 \gbuff_reg[9][30]  ( .D(n2477), .CK(clk), .RN(n1468), .Q(
        \gbuff[9][30] ) );
  DFFRX1 \gbuff_reg[9][29]  ( .D(n2478), .CK(clk), .RN(n1468), .Q(
        \gbuff[9][29] ) );
  DFFRX1 \gbuff_reg[9][28]  ( .D(n2479), .CK(clk), .RN(n1468), .Q(
        \gbuff[9][28] ) );
  DFFRX1 \gbuff_reg[9][27]  ( .D(n2480), .CK(clk), .RN(n1468), .Q(
        \gbuff[9][27] ) );
  DFFRX1 \gbuff_reg[9][26]  ( .D(n2481), .CK(clk), .RN(n1468), .Q(
        \gbuff[9][26] ) );
  DFFRX1 \gbuff_reg[9][25]  ( .D(n2482), .CK(clk), .RN(n1468), .Q(
        \gbuff[9][25] ) );
  DFFRX1 \gbuff_reg[9][24]  ( .D(n2483), .CK(clk), .RN(n1468), .Q(
        \gbuff[9][24] ) );
  DFFRX1 \gbuff_reg[9][23]  ( .D(n2484), .CK(clk), .RN(n1467), .Q(
        \gbuff[9][23] ) );
  DFFRX1 \gbuff_reg[9][22]  ( .D(n2485), .CK(clk), .RN(n1467), .Q(
        \gbuff[9][22] ) );
  DFFRX1 \gbuff_reg[9][21]  ( .D(n2486), .CK(clk), .RN(n1467), .Q(
        \gbuff[9][21] ) );
  DFFRX1 \gbuff_reg[9][20]  ( .D(n2487), .CK(clk), .RN(n1467), .Q(
        \gbuff[9][20] ) );
  DFFRX1 \gbuff_reg[9][19]  ( .D(n2488), .CK(clk), .RN(n1467), .Q(
        \gbuff[9][19] ) );
  DFFRX1 \gbuff_reg[9][18]  ( .D(n2489), .CK(clk), .RN(n1467), .Q(
        \gbuff[9][18] ) );
  DFFRX1 \gbuff_reg[9][17]  ( .D(n2490), .CK(clk), .RN(n1467), .Q(
        \gbuff[9][17] ) );
  DFFRX1 \gbuff_reg[9][16]  ( .D(n2491), .CK(clk), .RN(n1467), .Q(
        \gbuff[9][16] ) );
  DFFRX1 \gbuff_reg[9][15]  ( .D(n2492), .CK(clk), .RN(n1467), .Q(
        \gbuff[9][15] ) );
  DFFRX1 \gbuff_reg[9][14]  ( .D(n2493), .CK(clk), .RN(n1467), .Q(
        \gbuff[9][14] ) );
  DFFRX1 \gbuff_reg[9][13]  ( .D(n2494), .CK(clk), .RN(n1467), .Q(
        \gbuff[9][13] ) );
  DFFRX1 \gbuff_reg[9][12]  ( .D(n2495), .CK(clk), .RN(n1467), .Q(
        \gbuff[9][12] ) );
  DFFRX1 \gbuff_reg[9][11]  ( .D(n2496), .CK(clk), .RN(n1466), .Q(
        \gbuff[9][11] ) );
  DFFRX1 \gbuff_reg[9][10]  ( .D(n2497), .CK(clk), .RN(n1466), .Q(
        \gbuff[9][10] ) );
  DFFRX1 \gbuff_reg[9][9]  ( .D(n2498), .CK(clk), .RN(n1466), .Q(\gbuff[9][9] ) );
  DFFRX1 \gbuff_reg[9][8]  ( .D(n2499), .CK(clk), .RN(n1466), .Q(\gbuff[9][8] ) );
  DFFRX1 \gbuff_reg[9][7]  ( .D(n2500), .CK(clk), .RN(n1466), .Q(\gbuff[9][7] ) );
  DFFRX1 \gbuff_reg[9][6]  ( .D(n2501), .CK(clk), .RN(n1466), .Q(\gbuff[9][6] ) );
  DFFRX1 \gbuff_reg[9][5]  ( .D(n2502), .CK(clk), .RN(n1466), .Q(\gbuff[9][5] ) );
  DFFRX1 \gbuff_reg[9][4]  ( .D(n2503), .CK(clk), .RN(n1466), .Q(\gbuff[9][4] ) );
  DFFRX1 \gbuff_reg[9][3]  ( .D(n2504), .CK(clk), .RN(n1466), .Q(\gbuff[9][3] ) );
  DFFRX1 \gbuff_reg[9][2]  ( .D(n2505), .CK(clk), .RN(n1466), .Q(\gbuff[9][2] ) );
  DFFRX1 \gbuff_reg[9][1]  ( .D(n2506), .CK(clk), .RN(n1466), .Q(\gbuff[9][1] ) );
  DFFRX1 \gbuff_reg[9][0]  ( .D(n2507), .CK(clk), .RN(n1466), .Q(\gbuff[9][0] ) );
  DFFRX1 \gbuff_reg[5][31]  ( .D(n2604), .CK(clk), .RN(n1457), .Q(
        \gbuff[5][31] ) );
  DFFRX1 \gbuff_reg[5][30]  ( .D(n2605), .CK(clk), .RN(n1457), .Q(
        \gbuff[5][30] ) );
  DFFRX1 \gbuff_reg[5][29]  ( .D(n2606), .CK(clk), .RN(n1457), .Q(
        \gbuff[5][29] ) );
  DFFRX1 \gbuff_reg[5][28]  ( .D(n2607), .CK(clk), .RN(n1457), .Q(
        \gbuff[5][28] ) );
  DFFRX1 \gbuff_reg[5][27]  ( .D(n2608), .CK(clk), .RN(n1457), .Q(
        \gbuff[5][27] ) );
  DFFRX1 \gbuff_reg[5][26]  ( .D(n2609), .CK(clk), .RN(n1457), .Q(
        \gbuff[5][26] ) );
  DFFRX1 \gbuff_reg[5][25]  ( .D(n2610), .CK(clk), .RN(n1457), .Q(
        \gbuff[5][25] ) );
  DFFRX1 \gbuff_reg[5][24]  ( .D(n2611), .CK(clk), .RN(n1457), .Q(
        \gbuff[5][24] ) );
  DFFRX1 \gbuff_reg[5][23]  ( .D(n2612), .CK(clk), .RN(n1457), .Q(
        \gbuff[5][23] ) );
  DFFRX1 \gbuff_reg[5][22]  ( .D(n2613), .CK(clk), .RN(n1457), .Q(
        \gbuff[5][22] ) );
  DFFRX1 \gbuff_reg[5][21]  ( .D(n2614), .CK(clk), .RN(n1457), .Q(
        \gbuff[5][21] ) );
  DFFRX1 \gbuff_reg[5][20]  ( .D(n2615), .CK(clk), .RN(n1457), .Q(
        \gbuff[5][20] ) );
  DFFRX1 \gbuff_reg[5][19]  ( .D(n2616), .CK(clk), .RN(n1456), .Q(
        \gbuff[5][19] ) );
  DFFRX1 \gbuff_reg[5][18]  ( .D(n2617), .CK(clk), .RN(n1456), .Q(
        \gbuff[5][18] ) );
  DFFRX1 \gbuff_reg[5][17]  ( .D(n2618), .CK(clk), .RN(n1456), .Q(
        \gbuff[5][17] ) );
  DFFRX1 \gbuff_reg[5][16]  ( .D(n2619), .CK(clk), .RN(n1456), .Q(
        \gbuff[5][16] ) );
  DFFRX1 \gbuff_reg[5][15]  ( .D(n2620), .CK(clk), .RN(n1456), .Q(
        \gbuff[5][15] ) );
  DFFRX1 \gbuff_reg[5][14]  ( .D(n2621), .CK(clk), .RN(n1456), .Q(
        \gbuff[5][14] ) );
  DFFRX1 \gbuff_reg[5][13]  ( .D(n2622), .CK(clk), .RN(n1456), .Q(
        \gbuff[5][13] ) );
  DFFRX1 \gbuff_reg[5][12]  ( .D(n2623), .CK(clk), .RN(n1456), .Q(
        \gbuff[5][12] ) );
  DFFRX1 \gbuff_reg[5][11]  ( .D(n2624), .CK(clk), .RN(n1456), .Q(
        \gbuff[5][11] ) );
  DFFRX1 \gbuff_reg[5][10]  ( .D(n2625), .CK(clk), .RN(n1456), .Q(
        \gbuff[5][10] ) );
  DFFRX1 \gbuff_reg[5][9]  ( .D(n2626), .CK(clk), .RN(n1456), .Q(\gbuff[5][9] ) );
  DFFRX1 \gbuff_reg[5][8]  ( .D(n2627), .CK(clk), .RN(n1456), .Q(\gbuff[5][8] ) );
  DFFRX1 \gbuff_reg[5][7]  ( .D(n2628), .CK(clk), .RN(n1455), .Q(\gbuff[5][7] ) );
  DFFRX1 \gbuff_reg[5][6]  ( .D(n2629), .CK(clk), .RN(n1455), .Q(\gbuff[5][6] ) );
  DFFRX1 \gbuff_reg[5][5]  ( .D(n2630), .CK(clk), .RN(n1455), .Q(\gbuff[5][5] ) );
  DFFRX1 \gbuff_reg[5][4]  ( .D(n2631), .CK(clk), .RN(n1455), .Q(\gbuff[5][4] ) );
  DFFRX1 \gbuff_reg[5][3]  ( .D(n2632), .CK(clk), .RN(n1455), .Q(\gbuff[5][3] ) );
  DFFRX1 \gbuff_reg[5][2]  ( .D(n2633), .CK(clk), .RN(n1455), .Q(\gbuff[5][2] ) );
  DFFRX1 \gbuff_reg[5][1]  ( .D(n2634), .CK(clk), .RN(n1455), .Q(\gbuff[5][1] ) );
  DFFRX1 \gbuff_reg[5][0]  ( .D(n2635), .CK(clk), .RN(n1455), .Q(\gbuff[5][0] ) );
  DFFRX1 \gbuff_reg[1][31]  ( .D(n2732), .CK(clk), .RN(n1447), .Q(
        \gbuff[1][31] ) );
  DFFRX1 \gbuff_reg[1][30]  ( .D(n2733), .CK(clk), .RN(n1447), .Q(
        \gbuff[1][30] ) );
  DFFRX1 \gbuff_reg[1][29]  ( .D(n2734), .CK(clk), .RN(n1447), .Q(
        \gbuff[1][29] ) );
  DFFRX1 \gbuff_reg[1][28]  ( .D(n2735), .CK(clk), .RN(n1447), .Q(
        \gbuff[1][28] ) );
  DFFRX1 \gbuff_reg[1][27]  ( .D(n2736), .CK(clk), .RN(n1446), .Q(
        \gbuff[1][27] ) );
  DFFRX1 \gbuff_reg[1][26]  ( .D(n2737), .CK(clk), .RN(n1446), .Q(
        \gbuff[1][26] ) );
  DFFRX1 \gbuff_reg[1][25]  ( .D(n2738), .CK(clk), .RN(n1446), .Q(
        \gbuff[1][25] ) );
  DFFRX1 \gbuff_reg[1][24]  ( .D(n2739), .CK(clk), .RN(n1446), .Q(
        \gbuff[1][24] ) );
  DFFRX1 \gbuff_reg[1][23]  ( .D(n2740), .CK(clk), .RN(n1446), .Q(
        \gbuff[1][23] ) );
  DFFRX1 \gbuff_reg[1][22]  ( .D(n2741), .CK(clk), .RN(n1446), .Q(
        \gbuff[1][22] ) );
  DFFRX1 \gbuff_reg[1][21]  ( .D(n2742), .CK(clk), .RN(n1446), .Q(
        \gbuff[1][21] ) );
  DFFRX1 \gbuff_reg[1][20]  ( .D(n2743), .CK(clk), .RN(n1446), .Q(
        \gbuff[1][20] ) );
  DFFRX1 \gbuff_reg[1][19]  ( .D(n2744), .CK(clk), .RN(n1446), .Q(
        \gbuff[1][19] ) );
  DFFRX1 \gbuff_reg[1][18]  ( .D(n2745), .CK(clk), .RN(n1446), .Q(
        \gbuff[1][18] ) );
  DFFRX1 \gbuff_reg[1][17]  ( .D(n2746), .CK(clk), .RN(n1446), .Q(
        \gbuff[1][17] ) );
  DFFRX1 \gbuff_reg[1][16]  ( .D(n2747), .CK(clk), .RN(n1446), .Q(
        \gbuff[1][16] ) );
  DFFRX1 \gbuff_reg[1][15]  ( .D(n2748), .CK(clk), .RN(n1445), .Q(
        \gbuff[1][15] ) );
  DFFRX1 \gbuff_reg[1][14]  ( .D(n2749), .CK(clk), .RN(n1445), .Q(
        \gbuff[1][14] ) );
  DFFRX1 \gbuff_reg[1][13]  ( .D(n2750), .CK(clk), .RN(n1445), .Q(
        \gbuff[1][13] ) );
  DFFRX1 \gbuff_reg[1][12]  ( .D(n2751), .CK(clk), .RN(n1445), .Q(
        \gbuff[1][12] ) );
  DFFRX1 \gbuff_reg[1][11]  ( .D(n2752), .CK(clk), .RN(n1445), .Q(
        \gbuff[1][11] ) );
  DFFRX1 \gbuff_reg[1][10]  ( .D(n2753), .CK(clk), .RN(n1445), .Q(
        \gbuff[1][10] ) );
  DFFRX1 \gbuff_reg[1][9]  ( .D(n2754), .CK(clk), .RN(n1445), .Q(\gbuff[1][9] ) );
  DFFRX1 \gbuff_reg[1][8]  ( .D(n2755), .CK(clk), .RN(n1445), .Q(\gbuff[1][8] ) );
  DFFRX1 \gbuff_reg[1][7]  ( .D(n2756), .CK(clk), .RN(n1445), .Q(\gbuff[1][7] ) );
  DFFRX1 \gbuff_reg[1][6]  ( .D(n2757), .CK(clk), .RN(n1445), .Q(\gbuff[1][6] ) );
  DFFRX1 \gbuff_reg[1][5]  ( .D(n2758), .CK(clk), .RN(n1445), .Q(\gbuff[1][5] ) );
  DFFRX1 \gbuff_reg[1][4]  ( .D(n2759), .CK(clk), .RN(n1445), .Q(\gbuff[1][4] ) );
  DFFRX1 \gbuff_reg[1][3]  ( .D(n2760), .CK(clk), .RN(n1444), .Q(\gbuff[1][3] ) );
  DFFRX1 \gbuff_reg[1][2]  ( .D(n2761), .CK(clk), .RN(n1444), .Q(\gbuff[1][2] ) );
  DFFRX1 \gbuff_reg[1][1]  ( .D(n2762), .CK(clk), .RN(n1444), .Q(\gbuff[1][1] ) );
  DFFRX1 \gbuff_reg[1][0]  ( .D(n2763), .CK(clk), .RN(n1444), .Q(\gbuff[1][0] ) );
  DFFRX1 \gbuff_reg[31][31]  ( .D(n1772), .CK(clk), .RN(n1527), .Q(
        \gbuff[31][31] ) );
  DFFRX1 \gbuff_reg[31][30]  ( .D(n1773), .CK(clk), .RN(n1527), .Q(
        \gbuff[31][30] ) );
  DFFRX1 \gbuff_reg[31][29]  ( .D(n1774), .CK(clk), .RN(n1527), .Q(
        \gbuff[31][29] ) );
  DFFRX1 \gbuff_reg[31][28]  ( .D(n1775), .CK(clk), .RN(n1527), .Q(
        \gbuff[31][28] ) );
  DFFRX1 \gbuff_reg[31][27]  ( .D(n1776), .CK(clk), .RN(n1526), .Q(
        \gbuff[31][27] ) );
  DFFRX1 \gbuff_reg[31][26]  ( .D(n1777), .CK(clk), .RN(n1526), .Q(
        \gbuff[31][26] ) );
  DFFRX1 \gbuff_reg[31][25]  ( .D(n1778), .CK(clk), .RN(n1526), .Q(
        \gbuff[31][25] ) );
  DFFRX1 \gbuff_reg[31][24]  ( .D(n1779), .CK(clk), .RN(n1526), .Q(
        \gbuff[31][24] ) );
  DFFRX1 \gbuff_reg[31][23]  ( .D(n1780), .CK(clk), .RN(n1526), .Q(
        \gbuff[31][23] ) );
  DFFRX1 \gbuff_reg[31][22]  ( .D(n1781), .CK(clk), .RN(n1526), .Q(
        \gbuff[31][22] ) );
  DFFRX1 \gbuff_reg[31][21]  ( .D(n1782), .CK(clk), .RN(n1526), .Q(
        \gbuff[31][21] ) );
  DFFRX1 \gbuff_reg[31][20]  ( .D(n1783), .CK(clk), .RN(n1526), .Q(
        \gbuff[31][20] ) );
  DFFRX1 \gbuff_reg[31][19]  ( .D(n1784), .CK(clk), .RN(n1526), .Q(
        \gbuff[31][19] ) );
  DFFRX1 \gbuff_reg[31][18]  ( .D(n1785), .CK(clk), .RN(n1526), .Q(
        \gbuff[31][18] ) );
  DFFRX1 \gbuff_reg[31][17]  ( .D(n1786), .CK(clk), .RN(n1526), .Q(
        \gbuff[31][17] ) );
  DFFRX1 \gbuff_reg[31][16]  ( .D(n1787), .CK(clk), .RN(n1526), .Q(
        \gbuff[31][16] ) );
  DFFRX1 \gbuff_reg[31][15]  ( .D(n1788), .CK(clk), .RN(n1525), .Q(
        \gbuff[31][15] ) );
  DFFRX1 \gbuff_reg[31][14]  ( .D(n1789), .CK(clk), .RN(n1525), .Q(
        \gbuff[31][14] ) );
  DFFRX1 \gbuff_reg[31][13]  ( .D(n1790), .CK(clk), .RN(n1525), .Q(
        \gbuff[31][13] ) );
  DFFRX1 \gbuff_reg[31][12]  ( .D(n1791), .CK(clk), .RN(n1525), .Q(
        \gbuff[31][12] ) );
  DFFRX1 \gbuff_reg[31][11]  ( .D(n1792), .CK(clk), .RN(n1525), .Q(
        \gbuff[31][11] ) );
  DFFRX1 \gbuff_reg[31][10]  ( .D(n1793), .CK(clk), .RN(n1525), .Q(
        \gbuff[31][10] ) );
  DFFRX1 \gbuff_reg[31][9]  ( .D(n1794), .CK(clk), .RN(n1525), .Q(
        \gbuff[31][9] ) );
  DFFRX1 \gbuff_reg[31][8]  ( .D(n1795), .CK(clk), .RN(n1525), .Q(
        \gbuff[31][8] ) );
  DFFRX1 \gbuff_reg[31][7]  ( .D(n1796), .CK(clk), .RN(n1525), .Q(
        \gbuff[31][7] ) );
  DFFRX1 \gbuff_reg[31][6]  ( .D(n1797), .CK(clk), .RN(n1525), .Q(
        \gbuff[31][6] ) );
  DFFRX1 \gbuff_reg[31][5]  ( .D(n1798), .CK(clk), .RN(n1525), .Q(
        \gbuff[31][5] ) );
  DFFRX1 \gbuff_reg[31][4]  ( .D(n1799), .CK(clk), .RN(n1525), .Q(
        \gbuff[31][4] ) );
  DFFRX1 \gbuff_reg[31][3]  ( .D(n1800), .CK(clk), .RN(n1524), .Q(
        \gbuff[31][3] ) );
  DFFRX1 \gbuff_reg[31][2]  ( .D(n1801), .CK(clk), .RN(n1524), .Q(
        \gbuff[31][2] ) );
  DFFRX1 \gbuff_reg[31][1]  ( .D(n1802), .CK(clk), .RN(n1524), .Q(
        \gbuff[31][1] ) );
  DFFRX1 \gbuff_reg[31][0]  ( .D(n1803), .CK(clk), .RN(n1524), .Q(
        \gbuff[31][0] ) );
  DFFRX1 \gbuff_reg[27][31]  ( .D(n1900), .CK(clk), .RN(n1516), .Q(
        \gbuff[27][31] ) );
  DFFRX1 \gbuff_reg[27][30]  ( .D(n1901), .CK(clk), .RN(n1516), .Q(
        \gbuff[27][30] ) );
  DFFRX1 \gbuff_reg[27][29]  ( .D(n1902), .CK(clk), .RN(n1516), .Q(
        \gbuff[27][29] ) );
  DFFRX1 \gbuff_reg[27][28]  ( .D(n1903), .CK(clk), .RN(n1516), .Q(
        \gbuff[27][28] ) );
  DFFRX1 \gbuff_reg[27][27]  ( .D(n1904), .CK(clk), .RN(n1516), .Q(
        \gbuff[27][27] ) );
  DFFRX1 \gbuff_reg[27][26]  ( .D(n1905), .CK(clk), .RN(n1516), .Q(
        \gbuff[27][26] ) );
  DFFRX1 \gbuff_reg[27][25]  ( .D(n1906), .CK(clk), .RN(n1516), .Q(
        \gbuff[27][25] ) );
  DFFRX1 \gbuff_reg[27][24]  ( .D(n1907), .CK(clk), .RN(n1516), .Q(
        \gbuff[27][24] ) );
  DFFRX1 \gbuff_reg[27][23]  ( .D(n1908), .CK(clk), .RN(n1515), .Q(
        \gbuff[27][23] ) );
  DFFRX1 \gbuff_reg[27][22]  ( .D(n1909), .CK(clk), .RN(n1515), .Q(
        \gbuff[27][22] ) );
  DFFRX1 \gbuff_reg[27][21]  ( .D(n1910), .CK(clk), .RN(n1515), .Q(
        \gbuff[27][21] ) );
  DFFRX1 \gbuff_reg[27][20]  ( .D(n1911), .CK(clk), .RN(n1515), .Q(
        \gbuff[27][20] ) );
  DFFRX1 \gbuff_reg[27][19]  ( .D(n1912), .CK(clk), .RN(n1515), .Q(
        \gbuff[27][19] ) );
  DFFRX1 \gbuff_reg[27][18]  ( .D(n1913), .CK(clk), .RN(n1515), .Q(
        \gbuff[27][18] ) );
  DFFRX1 \gbuff_reg[27][17]  ( .D(n1914), .CK(clk), .RN(n1515), .Q(
        \gbuff[27][17] ) );
  DFFRX1 \gbuff_reg[27][16]  ( .D(n1915), .CK(clk), .RN(n1515), .Q(
        \gbuff[27][16] ) );
  DFFRX1 \gbuff_reg[27][15]  ( .D(n1916), .CK(clk), .RN(n1515), .Q(
        \gbuff[27][15] ) );
  DFFRX1 \gbuff_reg[27][14]  ( .D(n1917), .CK(clk), .RN(n1515), .Q(
        \gbuff[27][14] ) );
  DFFRX1 \gbuff_reg[27][13]  ( .D(n1918), .CK(clk), .RN(n1515), .Q(
        \gbuff[27][13] ) );
  DFFRX1 \gbuff_reg[27][12]  ( .D(n1919), .CK(clk), .RN(n1515), .Q(
        \gbuff[27][12] ) );
  DFFRX1 \gbuff_reg[27][11]  ( .D(n1920), .CK(clk), .RN(n1514), .Q(
        \gbuff[27][11] ) );
  DFFRX1 \gbuff_reg[27][10]  ( .D(n1921), .CK(clk), .RN(n1514), .Q(
        \gbuff[27][10] ) );
  DFFRX1 \gbuff_reg[27][9]  ( .D(n1922), .CK(clk), .RN(n1514), .Q(
        \gbuff[27][9] ) );
  DFFRX1 \gbuff_reg[27][8]  ( .D(n1923), .CK(clk), .RN(n1514), .Q(
        \gbuff[27][8] ) );
  DFFRX1 \gbuff_reg[27][7]  ( .D(n1924), .CK(clk), .RN(n1514), .Q(
        \gbuff[27][7] ) );
  DFFRX1 \gbuff_reg[27][6]  ( .D(n1925), .CK(clk), .RN(n1514), .Q(
        \gbuff[27][6] ) );
  DFFRX1 \gbuff_reg[27][5]  ( .D(n1926), .CK(clk), .RN(n1514), .Q(
        \gbuff[27][5] ) );
  DFFRX1 \gbuff_reg[27][4]  ( .D(n1927), .CK(clk), .RN(n1514), .Q(
        \gbuff[27][4] ) );
  DFFRX1 \gbuff_reg[27][3]  ( .D(n1928), .CK(clk), .RN(n1514), .Q(
        \gbuff[27][3] ) );
  DFFRX1 \gbuff_reg[27][2]  ( .D(n1929), .CK(clk), .RN(n1514), .Q(
        \gbuff[27][2] ) );
  DFFRX1 \gbuff_reg[27][1]  ( .D(n1930), .CK(clk), .RN(n1514), .Q(
        \gbuff[27][1] ) );
  DFFRX1 \gbuff_reg[27][0]  ( .D(n1931), .CK(clk), .RN(n1514), .Q(
        \gbuff[27][0] ) );
  DFFRX1 \gbuff_reg[23][31]  ( .D(n2028), .CK(clk), .RN(n1505), .Q(
        \gbuff[23][31] ) );
  DFFRX1 \gbuff_reg[23][30]  ( .D(n2029), .CK(clk), .RN(n1505), .Q(
        \gbuff[23][30] ) );
  DFFRX1 \gbuff_reg[23][29]  ( .D(n2030), .CK(clk), .RN(n1505), .Q(
        \gbuff[23][29] ) );
  DFFRX1 \gbuff_reg[23][28]  ( .D(n2031), .CK(clk), .RN(n1505), .Q(
        \gbuff[23][28] ) );
  DFFRX1 \gbuff_reg[23][27]  ( .D(n2032), .CK(clk), .RN(n1505), .Q(
        \gbuff[23][27] ) );
  DFFRX1 \gbuff_reg[23][26]  ( .D(n2033), .CK(clk), .RN(n1505), .Q(
        \gbuff[23][26] ) );
  DFFRX1 \gbuff_reg[23][25]  ( .D(n2034), .CK(clk), .RN(n1505), .Q(
        \gbuff[23][25] ) );
  DFFRX1 \gbuff_reg[23][24]  ( .D(n2035), .CK(clk), .RN(n1505), .Q(
        \gbuff[23][24] ) );
  DFFRX1 \gbuff_reg[23][23]  ( .D(n2036), .CK(clk), .RN(n1505), .Q(
        \gbuff[23][23] ) );
  DFFRX1 \gbuff_reg[23][22]  ( .D(n2037), .CK(clk), .RN(n1505), .Q(
        \gbuff[23][22] ) );
  DFFRX1 \gbuff_reg[23][21]  ( .D(n2038), .CK(clk), .RN(n1505), .Q(
        \gbuff[23][21] ) );
  DFFRX1 \gbuff_reg[23][20]  ( .D(n2039), .CK(clk), .RN(n1505), .Q(
        \gbuff[23][20] ) );
  DFFRX1 \gbuff_reg[23][19]  ( .D(n2040), .CK(clk), .RN(n1504), .Q(
        \gbuff[23][19] ) );
  DFFRX1 \gbuff_reg[23][18]  ( .D(n2041), .CK(clk), .RN(n1504), .Q(
        \gbuff[23][18] ) );
  DFFRX1 \gbuff_reg[23][17]  ( .D(n2042), .CK(clk), .RN(n1504), .Q(
        \gbuff[23][17] ) );
  DFFRX1 \gbuff_reg[23][16]  ( .D(n2043), .CK(clk), .RN(n1504), .Q(
        \gbuff[23][16] ) );
  DFFRX1 \gbuff_reg[23][15]  ( .D(n2044), .CK(clk), .RN(n1504), .Q(
        \gbuff[23][15] ) );
  DFFRX1 \gbuff_reg[23][14]  ( .D(n2045), .CK(clk), .RN(n1504), .Q(
        \gbuff[23][14] ) );
  DFFRX1 \gbuff_reg[23][13]  ( .D(n2046), .CK(clk), .RN(n1504), .Q(
        \gbuff[23][13] ) );
  DFFRX1 \gbuff_reg[23][12]  ( .D(n2047), .CK(clk), .RN(n1504), .Q(
        \gbuff[23][12] ) );
  DFFRX1 \gbuff_reg[23][11]  ( .D(n2048), .CK(clk), .RN(n1504), .Q(
        \gbuff[23][11] ) );
  DFFRX1 \gbuff_reg[23][10]  ( .D(n2049), .CK(clk), .RN(n1504), .Q(
        \gbuff[23][10] ) );
  DFFRX1 \gbuff_reg[23][9]  ( .D(n2050), .CK(clk), .RN(n1504), .Q(
        \gbuff[23][9] ) );
  DFFRX1 \gbuff_reg[23][8]  ( .D(n2051), .CK(clk), .RN(n1504), .Q(
        \gbuff[23][8] ) );
  DFFRX1 \gbuff_reg[23][7]  ( .D(n2052), .CK(clk), .RN(n1503), .Q(
        \gbuff[23][7] ) );
  DFFRX1 \gbuff_reg[23][6]  ( .D(n2053), .CK(clk), .RN(n1503), .Q(
        \gbuff[23][6] ) );
  DFFRX1 \gbuff_reg[23][5]  ( .D(n2054), .CK(clk), .RN(n1503), .Q(
        \gbuff[23][5] ) );
  DFFRX1 \gbuff_reg[23][4]  ( .D(n2055), .CK(clk), .RN(n1503), .Q(
        \gbuff[23][4] ) );
  DFFRX1 \gbuff_reg[23][3]  ( .D(n2056), .CK(clk), .RN(n1503), .Q(
        \gbuff[23][3] ) );
  DFFRX1 \gbuff_reg[23][2]  ( .D(n2057), .CK(clk), .RN(n1503), .Q(
        \gbuff[23][2] ) );
  DFFRX1 \gbuff_reg[23][1]  ( .D(n2058), .CK(clk), .RN(n1503), .Q(
        \gbuff[23][1] ) );
  DFFRX1 \gbuff_reg[23][0]  ( .D(n2059), .CK(clk), .RN(n1503), .Q(
        \gbuff[23][0] ) );
  DFFRX1 \gbuff_reg[19][31]  ( .D(n2156), .CK(clk), .RN(n1495), .Q(
        \gbuff[19][31] ) );
  DFFRX1 \gbuff_reg[19][30]  ( .D(n2157), .CK(clk), .RN(n1495), .Q(
        \gbuff[19][30] ) );
  DFFRX1 \gbuff_reg[19][29]  ( .D(n2158), .CK(clk), .RN(n1495), .Q(
        \gbuff[19][29] ) );
  DFFRX1 \gbuff_reg[19][28]  ( .D(n2159), .CK(clk), .RN(n1495), .Q(
        \gbuff[19][28] ) );
  DFFRX1 \gbuff_reg[19][27]  ( .D(n2160), .CK(clk), .RN(n1494), .Q(
        \gbuff[19][27] ) );
  DFFRX1 \gbuff_reg[19][26]  ( .D(n2161), .CK(clk), .RN(n1494), .Q(
        \gbuff[19][26] ) );
  DFFRX1 \gbuff_reg[19][25]  ( .D(n2162), .CK(clk), .RN(n1494), .Q(
        \gbuff[19][25] ) );
  DFFRX1 \gbuff_reg[19][24]  ( .D(n2163), .CK(clk), .RN(n1494), .Q(
        \gbuff[19][24] ) );
  DFFRX1 \gbuff_reg[19][23]  ( .D(n2164), .CK(clk), .RN(n1494), .Q(
        \gbuff[19][23] ) );
  DFFRX1 \gbuff_reg[19][22]  ( .D(n2165), .CK(clk), .RN(n1494), .Q(
        \gbuff[19][22] ) );
  DFFRX1 \gbuff_reg[19][21]  ( .D(n2166), .CK(clk), .RN(n1494), .Q(
        \gbuff[19][21] ) );
  DFFRX1 \gbuff_reg[19][20]  ( .D(n2167), .CK(clk), .RN(n1494), .Q(
        \gbuff[19][20] ) );
  DFFRX1 \gbuff_reg[19][19]  ( .D(n2168), .CK(clk), .RN(n1494), .Q(
        \gbuff[19][19] ) );
  DFFRX1 \gbuff_reg[19][18]  ( .D(n2169), .CK(clk), .RN(n1494), .Q(
        \gbuff[19][18] ) );
  DFFRX1 \gbuff_reg[19][17]  ( .D(n2170), .CK(clk), .RN(n1494), .Q(
        \gbuff[19][17] ) );
  DFFRX1 \gbuff_reg[19][16]  ( .D(n2171), .CK(clk), .RN(n1494), .Q(
        \gbuff[19][16] ) );
  DFFRX1 \gbuff_reg[19][15]  ( .D(n2172), .CK(clk), .RN(n1493), .Q(
        \gbuff[19][15] ) );
  DFFRX1 \gbuff_reg[19][14]  ( .D(n2173), .CK(clk), .RN(n1493), .Q(
        \gbuff[19][14] ) );
  DFFRX1 \gbuff_reg[19][13]  ( .D(n2174), .CK(clk), .RN(n1493), .Q(
        \gbuff[19][13] ) );
  DFFRX1 \gbuff_reg[19][12]  ( .D(n2175), .CK(clk), .RN(n1493), .Q(
        \gbuff[19][12] ) );
  DFFRX1 \gbuff_reg[19][11]  ( .D(n2176), .CK(clk), .RN(n1493), .Q(
        \gbuff[19][11] ) );
  DFFRX1 \gbuff_reg[19][10]  ( .D(n2177), .CK(clk), .RN(n1493), .Q(
        \gbuff[19][10] ) );
  DFFRX1 \gbuff_reg[19][9]  ( .D(n2178), .CK(clk), .RN(n1493), .Q(
        \gbuff[19][9] ) );
  DFFRX1 \gbuff_reg[19][8]  ( .D(n2179), .CK(clk), .RN(n1493), .Q(
        \gbuff[19][8] ) );
  DFFRX1 \gbuff_reg[19][7]  ( .D(n2180), .CK(clk), .RN(n1493), .Q(
        \gbuff[19][7] ) );
  DFFRX1 \gbuff_reg[19][6]  ( .D(n2181), .CK(clk), .RN(n1493), .Q(
        \gbuff[19][6] ) );
  DFFRX1 \gbuff_reg[19][5]  ( .D(n2182), .CK(clk), .RN(n1493), .Q(
        \gbuff[19][5] ) );
  DFFRX1 \gbuff_reg[19][4]  ( .D(n2183), .CK(clk), .RN(n1493), .Q(
        \gbuff[19][4] ) );
  DFFRX1 \gbuff_reg[19][3]  ( .D(n2184), .CK(clk), .RN(n1492), .Q(
        \gbuff[19][3] ) );
  DFFRX1 \gbuff_reg[19][2]  ( .D(n2185), .CK(clk), .RN(n1492), .Q(
        \gbuff[19][2] ) );
  DFFRX1 \gbuff_reg[19][1]  ( .D(n2186), .CK(clk), .RN(n1492), .Q(
        \gbuff[19][1] ) );
  DFFRX1 \gbuff_reg[19][0]  ( .D(n2187), .CK(clk), .RN(n1492), .Q(
        \gbuff[19][0] ) );
  DFFRX1 \gbuff_reg[15][31]  ( .D(n2284), .CK(clk), .RN(n1484), .Q(
        \gbuff[15][31] ) );
  DFFRX1 \gbuff_reg[15][30]  ( .D(n2285), .CK(clk), .RN(n1484), .Q(
        \gbuff[15][30] ) );
  DFFRX1 \gbuff_reg[15][29]  ( .D(n2286), .CK(clk), .RN(n1484), .Q(
        \gbuff[15][29] ) );
  DFFRX1 \gbuff_reg[15][28]  ( .D(n2287), .CK(clk), .RN(n1484), .Q(
        \gbuff[15][28] ) );
  DFFRX1 \gbuff_reg[15][27]  ( .D(n2288), .CK(clk), .RN(n1484), .Q(
        \gbuff[15][27] ) );
  DFFRX1 \gbuff_reg[15][26]  ( .D(n2289), .CK(clk), .RN(n1484), .Q(
        \gbuff[15][26] ) );
  DFFRX1 \gbuff_reg[15][25]  ( .D(n2290), .CK(clk), .RN(n1484), .Q(
        \gbuff[15][25] ) );
  DFFRX1 \gbuff_reg[15][24]  ( .D(n2291), .CK(clk), .RN(n1484), .Q(
        \gbuff[15][24] ) );
  DFFRX1 \gbuff_reg[15][23]  ( .D(n2292), .CK(clk), .RN(n1483), .Q(
        \gbuff[15][23] ) );
  DFFRX1 \gbuff_reg[15][22]  ( .D(n2293), .CK(clk), .RN(n1483), .Q(
        \gbuff[15][22] ) );
  DFFRX1 \gbuff_reg[15][21]  ( .D(n2294), .CK(clk), .RN(n1483), .Q(
        \gbuff[15][21] ) );
  DFFRX1 \gbuff_reg[15][20]  ( .D(n2295), .CK(clk), .RN(n1483), .Q(
        \gbuff[15][20] ) );
  DFFRX1 \gbuff_reg[15][19]  ( .D(n2296), .CK(clk), .RN(n1483), .Q(
        \gbuff[15][19] ) );
  DFFRX1 \gbuff_reg[15][18]  ( .D(n2297), .CK(clk), .RN(n1483), .Q(
        \gbuff[15][18] ) );
  DFFRX1 \gbuff_reg[15][17]  ( .D(n2298), .CK(clk), .RN(n1483), .Q(
        \gbuff[15][17] ) );
  DFFRX1 \gbuff_reg[15][16]  ( .D(n2299), .CK(clk), .RN(n1483), .Q(
        \gbuff[15][16] ) );
  DFFRX1 \gbuff_reg[15][15]  ( .D(n2300), .CK(clk), .RN(n1483), .Q(
        \gbuff[15][15] ) );
  DFFRX1 \gbuff_reg[15][14]  ( .D(n2301), .CK(clk), .RN(n1483), .Q(
        \gbuff[15][14] ) );
  DFFRX1 \gbuff_reg[15][13]  ( .D(n2302), .CK(clk), .RN(n1483), .Q(
        \gbuff[15][13] ) );
  DFFRX1 \gbuff_reg[15][12]  ( .D(n2303), .CK(clk), .RN(n1483), .Q(
        \gbuff[15][12] ) );
  DFFRX1 \gbuff_reg[15][11]  ( .D(n2304), .CK(clk), .RN(n1482), .Q(
        \gbuff[15][11] ) );
  DFFRX1 \gbuff_reg[15][10]  ( .D(n2305), .CK(clk), .RN(n1482), .Q(
        \gbuff[15][10] ) );
  DFFRX1 \gbuff_reg[15][9]  ( .D(n2306), .CK(clk), .RN(n1482), .Q(
        \gbuff[15][9] ) );
  DFFRX1 \gbuff_reg[15][8]  ( .D(n2307), .CK(clk), .RN(n1482), .Q(
        \gbuff[15][8] ) );
  DFFRX1 \gbuff_reg[15][7]  ( .D(n2308), .CK(clk), .RN(n1482), .Q(
        \gbuff[15][7] ) );
  DFFRX1 \gbuff_reg[15][6]  ( .D(n2309), .CK(clk), .RN(n1482), .Q(
        \gbuff[15][6] ) );
  DFFRX1 \gbuff_reg[15][5]  ( .D(n2310), .CK(clk), .RN(n1482), .Q(
        \gbuff[15][5] ) );
  DFFRX1 \gbuff_reg[15][4]  ( .D(n2311), .CK(clk), .RN(n1482), .Q(
        \gbuff[15][4] ) );
  DFFRX1 \gbuff_reg[15][3]  ( .D(n2312), .CK(clk), .RN(n1482), .Q(
        \gbuff[15][3] ) );
  DFFRX1 \gbuff_reg[15][2]  ( .D(n2313), .CK(clk), .RN(n1482), .Q(
        \gbuff[15][2] ) );
  DFFRX1 \gbuff_reg[15][1]  ( .D(n2314), .CK(clk), .RN(n1482), .Q(
        \gbuff[15][1] ) );
  DFFRX1 \gbuff_reg[15][0]  ( .D(n2315), .CK(clk), .RN(n1482), .Q(
        \gbuff[15][0] ) );
  DFFRX1 \gbuff_reg[11][31]  ( .D(n2412), .CK(clk), .RN(n1473), .Q(
        \gbuff[11][31] ) );
  DFFRX1 \gbuff_reg[11][30]  ( .D(n2413), .CK(clk), .RN(n1473), .Q(
        \gbuff[11][30] ) );
  DFFRX1 \gbuff_reg[11][29]  ( .D(n2414), .CK(clk), .RN(n1473), .Q(
        \gbuff[11][29] ) );
  DFFRX1 \gbuff_reg[11][28]  ( .D(n2415), .CK(clk), .RN(n1473), .Q(
        \gbuff[11][28] ) );
  DFFRX1 \gbuff_reg[11][27]  ( .D(n2416), .CK(clk), .RN(n1473), .Q(
        \gbuff[11][27] ) );
  DFFRX1 \gbuff_reg[11][26]  ( .D(n2417), .CK(clk), .RN(n1473), .Q(
        \gbuff[11][26] ) );
  DFFRX1 \gbuff_reg[11][25]  ( .D(n2418), .CK(clk), .RN(n1473), .Q(
        \gbuff[11][25] ) );
  DFFRX1 \gbuff_reg[11][24]  ( .D(n2419), .CK(clk), .RN(n1473), .Q(
        \gbuff[11][24] ) );
  DFFRX1 \gbuff_reg[11][23]  ( .D(n2420), .CK(clk), .RN(n1473), .Q(
        \gbuff[11][23] ) );
  DFFRX1 \gbuff_reg[11][22]  ( .D(n2421), .CK(clk), .RN(n1473), .Q(
        \gbuff[11][22] ) );
  DFFRX1 \gbuff_reg[11][21]  ( .D(n2422), .CK(clk), .RN(n1473), .Q(
        \gbuff[11][21] ) );
  DFFRX1 \gbuff_reg[11][20]  ( .D(n2423), .CK(clk), .RN(n1473), .Q(
        \gbuff[11][20] ) );
  DFFRX1 \gbuff_reg[11][19]  ( .D(n2424), .CK(clk), .RN(n1472), .Q(
        \gbuff[11][19] ) );
  DFFRX1 \gbuff_reg[11][18]  ( .D(n2425), .CK(clk), .RN(n1472), .Q(
        \gbuff[11][18] ) );
  DFFRX1 \gbuff_reg[11][17]  ( .D(n2426), .CK(clk), .RN(n1472), .Q(
        \gbuff[11][17] ) );
  DFFRX1 \gbuff_reg[11][16]  ( .D(n2427), .CK(clk), .RN(n1472), .Q(
        \gbuff[11][16] ) );
  DFFRX1 \gbuff_reg[11][15]  ( .D(n2428), .CK(clk), .RN(n1472), .Q(
        \gbuff[11][15] ) );
  DFFRX1 \gbuff_reg[11][14]  ( .D(n2429), .CK(clk), .RN(n1472), .Q(
        \gbuff[11][14] ) );
  DFFRX1 \gbuff_reg[11][13]  ( .D(n2430), .CK(clk), .RN(n1472), .Q(
        \gbuff[11][13] ) );
  DFFRX1 \gbuff_reg[11][12]  ( .D(n2431), .CK(clk), .RN(n1472), .Q(
        \gbuff[11][12] ) );
  DFFRX1 \gbuff_reg[11][11]  ( .D(n2432), .CK(clk), .RN(n1472), .Q(
        \gbuff[11][11] ) );
  DFFRX1 \gbuff_reg[11][10]  ( .D(n2433), .CK(clk), .RN(n1472), .Q(
        \gbuff[11][10] ) );
  DFFRX1 \gbuff_reg[11][9]  ( .D(n2434), .CK(clk), .RN(n1472), .Q(
        \gbuff[11][9] ) );
  DFFRX1 \gbuff_reg[11][8]  ( .D(n2435), .CK(clk), .RN(n1472), .Q(
        \gbuff[11][8] ) );
  DFFRX1 \gbuff_reg[11][7]  ( .D(n2436), .CK(clk), .RN(n1471), .Q(
        \gbuff[11][7] ) );
  DFFRX1 \gbuff_reg[11][6]  ( .D(n2437), .CK(clk), .RN(n1471), .Q(
        \gbuff[11][6] ) );
  DFFRX1 \gbuff_reg[11][5]  ( .D(n2438), .CK(clk), .RN(n1471), .Q(
        \gbuff[11][5] ) );
  DFFRX1 \gbuff_reg[11][4]  ( .D(n2439), .CK(clk), .RN(n1471), .Q(
        \gbuff[11][4] ) );
  DFFRX1 \gbuff_reg[11][3]  ( .D(n2440), .CK(clk), .RN(n1471), .Q(
        \gbuff[11][3] ) );
  DFFRX1 \gbuff_reg[11][2]  ( .D(n2441), .CK(clk), .RN(n1471), .Q(
        \gbuff[11][2] ) );
  DFFRX1 \gbuff_reg[11][1]  ( .D(n2442), .CK(clk), .RN(n1471), .Q(
        \gbuff[11][1] ) );
  DFFRX1 \gbuff_reg[11][0]  ( .D(n2443), .CK(clk), .RN(n1471), .Q(
        \gbuff[11][0] ) );
  DFFRX1 \gbuff_reg[7][31]  ( .D(n2540), .CK(clk), .RN(n1463), .Q(
        \gbuff[7][31] ) );
  DFFRX1 \gbuff_reg[7][30]  ( .D(n2541), .CK(clk), .RN(n1463), .Q(
        \gbuff[7][30] ) );
  DFFRX1 \gbuff_reg[7][29]  ( .D(n2542), .CK(clk), .RN(n1463), .Q(
        \gbuff[7][29] ) );
  DFFRX1 \gbuff_reg[7][28]  ( .D(n2543), .CK(clk), .RN(n1463), .Q(
        \gbuff[7][28] ) );
  DFFRX1 \gbuff_reg[7][27]  ( .D(n2544), .CK(clk), .RN(n1462), .Q(
        \gbuff[7][27] ) );
  DFFRX1 \gbuff_reg[7][26]  ( .D(n2545), .CK(clk), .RN(n1462), .Q(
        \gbuff[7][26] ) );
  DFFRX1 \gbuff_reg[7][25]  ( .D(n2546), .CK(clk), .RN(n1462), .Q(
        \gbuff[7][25] ) );
  DFFRX1 \gbuff_reg[7][24]  ( .D(n2547), .CK(clk), .RN(n1462), .Q(
        \gbuff[7][24] ) );
  DFFRX1 \gbuff_reg[7][23]  ( .D(n2548), .CK(clk), .RN(n1462), .Q(
        \gbuff[7][23] ) );
  DFFRX1 \gbuff_reg[7][22]  ( .D(n2549), .CK(clk), .RN(n1462), .Q(
        \gbuff[7][22] ) );
  DFFRX1 \gbuff_reg[7][21]  ( .D(n2550), .CK(clk), .RN(n1462), .Q(
        \gbuff[7][21] ) );
  DFFRX1 \gbuff_reg[7][20]  ( .D(n2551), .CK(clk), .RN(n1462), .Q(
        \gbuff[7][20] ) );
  DFFRX1 \gbuff_reg[7][19]  ( .D(n2552), .CK(clk), .RN(n1462), .Q(
        \gbuff[7][19] ) );
  DFFRX1 \gbuff_reg[7][18]  ( .D(n2553), .CK(clk), .RN(n1462), .Q(
        \gbuff[7][18] ) );
  DFFRX1 \gbuff_reg[7][17]  ( .D(n2554), .CK(clk), .RN(n1462), .Q(
        \gbuff[7][17] ) );
  DFFRX1 \gbuff_reg[7][16]  ( .D(n2555), .CK(clk), .RN(n1462), .Q(
        \gbuff[7][16] ) );
  DFFRX1 \gbuff_reg[7][15]  ( .D(n2556), .CK(clk), .RN(n1461), .Q(
        \gbuff[7][15] ) );
  DFFRX1 \gbuff_reg[7][14]  ( .D(n2557), .CK(clk), .RN(n1461), .Q(
        \gbuff[7][14] ) );
  DFFRX1 \gbuff_reg[7][13]  ( .D(n2558), .CK(clk), .RN(n1461), .Q(
        \gbuff[7][13] ) );
  DFFRX1 \gbuff_reg[7][12]  ( .D(n2559), .CK(clk), .RN(n1461), .Q(
        \gbuff[7][12] ) );
  DFFRX1 \gbuff_reg[7][11]  ( .D(n2560), .CK(clk), .RN(n1461), .Q(
        \gbuff[7][11] ) );
  DFFRX1 \gbuff_reg[7][10]  ( .D(n2561), .CK(clk), .RN(n1461), .Q(
        \gbuff[7][10] ) );
  DFFRX1 \gbuff_reg[7][9]  ( .D(n2562), .CK(clk), .RN(n1461), .Q(\gbuff[7][9] ) );
  DFFRX1 \gbuff_reg[7][8]  ( .D(n2563), .CK(clk), .RN(n1461), .Q(\gbuff[7][8] ) );
  DFFRX1 \gbuff_reg[7][7]  ( .D(n2564), .CK(clk), .RN(n1461), .Q(\gbuff[7][7] ) );
  DFFRX1 \gbuff_reg[7][6]  ( .D(n2565), .CK(clk), .RN(n1461), .Q(\gbuff[7][6] ) );
  DFFRX1 \gbuff_reg[7][5]  ( .D(n2566), .CK(clk), .RN(n1461), .Q(\gbuff[7][5] ) );
  DFFRX1 \gbuff_reg[7][4]  ( .D(n2567), .CK(clk), .RN(n1461), .Q(\gbuff[7][4] ) );
  DFFRX1 \gbuff_reg[7][3]  ( .D(n2568), .CK(clk), .RN(n1460), .Q(\gbuff[7][3] ) );
  DFFRX1 \gbuff_reg[7][2]  ( .D(n2569), .CK(clk), .RN(n1460), .Q(\gbuff[7][2] ) );
  DFFRX1 \gbuff_reg[7][1]  ( .D(n2570), .CK(clk), .RN(n1460), .Q(\gbuff[7][1] ) );
  DFFRX1 \gbuff_reg[7][0]  ( .D(n2571), .CK(clk), .RN(n1460), .Q(\gbuff[7][0] ) );
  DFFRX1 \gbuff_reg[3][31]  ( .D(n2668), .CK(clk), .RN(n1452), .Q(
        \gbuff[3][31] ) );
  DFFRX1 \gbuff_reg[3][30]  ( .D(n2669), .CK(clk), .RN(n1452), .Q(
        \gbuff[3][30] ) );
  DFFRX1 \gbuff_reg[3][29]  ( .D(n2670), .CK(clk), .RN(n1452), .Q(
        \gbuff[3][29] ) );
  DFFRX1 \gbuff_reg[3][28]  ( .D(n2671), .CK(clk), .RN(n1452), .Q(
        \gbuff[3][28] ) );
  DFFRX1 \gbuff_reg[3][27]  ( .D(n2672), .CK(clk), .RN(n1452), .Q(
        \gbuff[3][27] ) );
  DFFRX1 \gbuff_reg[3][26]  ( .D(n2673), .CK(clk), .RN(n1452), .Q(
        \gbuff[3][26] ) );
  DFFRX1 \gbuff_reg[3][25]  ( .D(n2674), .CK(clk), .RN(n1452), .Q(
        \gbuff[3][25] ) );
  DFFRX1 \gbuff_reg[3][24]  ( .D(n2675), .CK(clk), .RN(n1452), .Q(
        \gbuff[3][24] ) );
  DFFRX1 \gbuff_reg[3][23]  ( .D(n2676), .CK(clk), .RN(n1451), .Q(
        \gbuff[3][23] ) );
  DFFRX1 \gbuff_reg[3][22]  ( .D(n2677), .CK(clk), .RN(n1451), .Q(
        \gbuff[3][22] ) );
  DFFRX1 \gbuff_reg[3][21]  ( .D(n2678), .CK(clk), .RN(n1451), .Q(
        \gbuff[3][21] ) );
  DFFRX1 \gbuff_reg[3][20]  ( .D(n2679), .CK(clk), .RN(n1451), .Q(
        \gbuff[3][20] ) );
  DFFRX1 \gbuff_reg[3][19]  ( .D(n2680), .CK(clk), .RN(n1451), .Q(
        \gbuff[3][19] ) );
  DFFRX1 \gbuff_reg[3][18]  ( .D(n2681), .CK(clk), .RN(n1451), .Q(
        \gbuff[3][18] ) );
  DFFRX1 \gbuff_reg[3][17]  ( .D(n2682), .CK(clk), .RN(n1451), .Q(
        \gbuff[3][17] ) );
  DFFRX1 \gbuff_reg[3][16]  ( .D(n2683), .CK(clk), .RN(n1451), .Q(
        \gbuff[3][16] ) );
  DFFRX1 \gbuff_reg[3][15]  ( .D(n2684), .CK(clk), .RN(n1451), .Q(
        \gbuff[3][15] ) );
  DFFRX1 \gbuff_reg[3][14]  ( .D(n2685), .CK(clk), .RN(n1451), .Q(
        \gbuff[3][14] ) );
  DFFRX1 \gbuff_reg[3][13]  ( .D(n2686), .CK(clk), .RN(n1451), .Q(
        \gbuff[3][13] ) );
  DFFRX1 \gbuff_reg[3][12]  ( .D(n2687), .CK(clk), .RN(n1451), .Q(
        \gbuff[3][12] ) );
  DFFRX1 \gbuff_reg[3][11]  ( .D(n2688), .CK(clk), .RN(n1450), .Q(
        \gbuff[3][11] ) );
  DFFRX1 \gbuff_reg[3][10]  ( .D(n2689), .CK(clk), .RN(n1450), .Q(
        \gbuff[3][10] ) );
  DFFRX1 \gbuff_reg[3][9]  ( .D(n2690), .CK(clk), .RN(n1450), .Q(\gbuff[3][9] ) );
  DFFRX1 \gbuff_reg[3][8]  ( .D(n2691), .CK(clk), .RN(n1450), .Q(\gbuff[3][8] ) );
  DFFRX1 \gbuff_reg[3][7]  ( .D(n2692), .CK(clk), .RN(n1450), .Q(\gbuff[3][7] ) );
  DFFRX1 \gbuff_reg[3][6]  ( .D(n2693), .CK(clk), .RN(n1450), .Q(\gbuff[3][6] ) );
  DFFRX1 \gbuff_reg[3][5]  ( .D(n2694), .CK(clk), .RN(n1450), .Q(\gbuff[3][5] ) );
  DFFRX1 \gbuff_reg[3][4]  ( .D(n2695), .CK(clk), .RN(n1450), .Q(\gbuff[3][4] ) );
  DFFRX1 \gbuff_reg[3][3]  ( .D(n2696), .CK(clk), .RN(n1450), .Q(\gbuff[3][3] ) );
  DFFRX1 \gbuff_reg[3][2]  ( .D(n2697), .CK(clk), .RN(n1450), .Q(\gbuff[3][2] ) );
  DFFRX1 \gbuff_reg[3][1]  ( .D(n2698), .CK(clk), .RN(n1450), .Q(\gbuff[3][1] ) );
  DFFRX1 \gbuff_reg[3][0]  ( .D(n2699), .CK(clk), .RN(n1450), .Q(\gbuff[3][0] ) );
  DFFRX1 \gbuff_reg[28][31]  ( .D(n1868), .CK(clk), .RN(n1519), .Q(
        \gbuff[28][31] ) );
  DFFRX1 \gbuff_reg[28][30]  ( .D(n1869), .CK(clk), .RN(n1519), .Q(
        \gbuff[28][30] ) );
  DFFRX1 \gbuff_reg[28][29]  ( .D(n1870), .CK(clk), .RN(n1519), .Q(
        \gbuff[28][29] ) );
  DFFRX1 \gbuff_reg[28][28]  ( .D(n1871), .CK(clk), .RN(n1519), .Q(
        \gbuff[28][28] ) );
  DFFRX1 \gbuff_reg[28][27]  ( .D(n1872), .CK(clk), .RN(n1518), .Q(
        \gbuff[28][27] ) );
  DFFRX1 \gbuff_reg[28][26]  ( .D(n1873), .CK(clk), .RN(n1518), .Q(
        \gbuff[28][26] ) );
  DFFRX1 \gbuff_reg[28][25]  ( .D(n1874), .CK(clk), .RN(n1518), .Q(
        \gbuff[28][25] ) );
  DFFRX1 \gbuff_reg[28][24]  ( .D(n1875), .CK(clk), .RN(n1518), .Q(
        \gbuff[28][24] ) );
  DFFRX1 \gbuff_reg[28][23]  ( .D(n1876), .CK(clk), .RN(n1518), .Q(
        \gbuff[28][23] ) );
  DFFRX1 \gbuff_reg[28][22]  ( .D(n1877), .CK(clk), .RN(n1518), .Q(
        \gbuff[28][22] ) );
  DFFRX1 \gbuff_reg[28][21]  ( .D(n1878), .CK(clk), .RN(n1518), .Q(
        \gbuff[28][21] ) );
  DFFRX1 \gbuff_reg[28][20]  ( .D(n1879), .CK(clk), .RN(n1518), .Q(
        \gbuff[28][20] ) );
  DFFRX1 \gbuff_reg[28][19]  ( .D(n1880), .CK(clk), .RN(n1518), .Q(
        \gbuff[28][19] ) );
  DFFRX1 \gbuff_reg[28][18]  ( .D(n1881), .CK(clk), .RN(n1518), .Q(
        \gbuff[28][18] ) );
  DFFRX1 \gbuff_reg[28][17]  ( .D(n1882), .CK(clk), .RN(n1518), .Q(
        \gbuff[28][17] ) );
  DFFRX1 \gbuff_reg[28][16]  ( .D(n1883), .CK(clk), .RN(n1518), .Q(
        \gbuff[28][16] ) );
  DFFRX1 \gbuff_reg[28][15]  ( .D(n1884), .CK(clk), .RN(n1517), .Q(
        \gbuff[28][15] ) );
  DFFRX1 \gbuff_reg[28][14]  ( .D(n1885), .CK(clk), .RN(n1517), .Q(
        \gbuff[28][14] ) );
  DFFRX1 \gbuff_reg[28][13]  ( .D(n1886), .CK(clk), .RN(n1517), .Q(
        \gbuff[28][13] ) );
  DFFRX1 \gbuff_reg[28][12]  ( .D(n1887), .CK(clk), .RN(n1517), .Q(
        \gbuff[28][12] ) );
  DFFRX1 \gbuff_reg[28][11]  ( .D(n1888), .CK(clk), .RN(n1517), .Q(
        \gbuff[28][11] ) );
  DFFRX1 \gbuff_reg[28][10]  ( .D(n1889), .CK(clk), .RN(n1517), .Q(
        \gbuff[28][10] ) );
  DFFRX1 \gbuff_reg[28][9]  ( .D(n1890), .CK(clk), .RN(n1517), .Q(
        \gbuff[28][9] ) );
  DFFRX1 \gbuff_reg[28][8]  ( .D(n1891), .CK(clk), .RN(n1517), .Q(
        \gbuff[28][8] ) );
  DFFRX1 \gbuff_reg[28][7]  ( .D(n1892), .CK(clk), .RN(n1517), .Q(
        \gbuff[28][7] ) );
  DFFRX1 \gbuff_reg[28][6]  ( .D(n1893), .CK(clk), .RN(n1517), .Q(
        \gbuff[28][6] ) );
  DFFRX1 \gbuff_reg[28][5]  ( .D(n1894), .CK(clk), .RN(n1517), .Q(
        \gbuff[28][5] ) );
  DFFRX1 \gbuff_reg[28][4]  ( .D(n1895), .CK(clk), .RN(n1517), .Q(
        \gbuff[28][4] ) );
  DFFRX1 \gbuff_reg[28][3]  ( .D(n1896), .CK(clk), .RN(n1516), .Q(
        \gbuff[28][3] ) );
  DFFRX1 \gbuff_reg[28][2]  ( .D(n1897), .CK(clk), .RN(n1516), .Q(
        \gbuff[28][2] ) );
  DFFRX1 \gbuff_reg[28][1]  ( .D(n1898), .CK(clk), .RN(n1516), .Q(
        \gbuff[28][1] ) );
  DFFRX1 \gbuff_reg[28][0]  ( .D(n1899), .CK(clk), .RN(n1516), .Q(
        \gbuff[28][0] ) );
  DFFRX1 \gbuff_reg[24][31]  ( .D(n1996), .CK(clk), .RN(n1508), .Q(
        \gbuff[24][31] ) );
  DFFRX1 \gbuff_reg[24][30]  ( .D(n1997), .CK(clk), .RN(n1508), .Q(
        \gbuff[24][30] ) );
  DFFRX1 \gbuff_reg[24][29]  ( .D(n1998), .CK(clk), .RN(n1508), .Q(
        \gbuff[24][29] ) );
  DFFRX1 \gbuff_reg[24][28]  ( .D(n1999), .CK(clk), .RN(n1508), .Q(
        \gbuff[24][28] ) );
  DFFRX1 \gbuff_reg[24][27]  ( .D(n2000), .CK(clk), .RN(n1508), .Q(
        \gbuff[24][27] ) );
  DFFRX1 \gbuff_reg[24][26]  ( .D(n2001), .CK(clk), .RN(n1508), .Q(
        \gbuff[24][26] ) );
  DFFRX1 \gbuff_reg[24][25]  ( .D(n2002), .CK(clk), .RN(n1508), .Q(
        \gbuff[24][25] ) );
  DFFRX1 \gbuff_reg[24][24]  ( .D(n2003), .CK(clk), .RN(n1508), .Q(
        \gbuff[24][24] ) );
  DFFRX1 \gbuff_reg[24][23]  ( .D(n2004), .CK(clk), .RN(n1507), .Q(
        \gbuff[24][23] ) );
  DFFRX1 \gbuff_reg[24][22]  ( .D(n2005), .CK(clk), .RN(n1507), .Q(
        \gbuff[24][22] ) );
  DFFRX1 \gbuff_reg[24][21]  ( .D(n2006), .CK(clk), .RN(n1507), .Q(
        \gbuff[24][21] ) );
  DFFRX1 \gbuff_reg[24][20]  ( .D(n2007), .CK(clk), .RN(n1507), .Q(
        \gbuff[24][20] ) );
  DFFRX1 \gbuff_reg[24][19]  ( .D(n2008), .CK(clk), .RN(n1507), .Q(
        \gbuff[24][19] ) );
  DFFRX1 \gbuff_reg[24][18]  ( .D(n2009), .CK(clk), .RN(n1507), .Q(
        \gbuff[24][18] ) );
  DFFRX1 \gbuff_reg[24][17]  ( .D(n2010), .CK(clk), .RN(n1507), .Q(
        \gbuff[24][17] ) );
  DFFRX1 \gbuff_reg[24][16]  ( .D(n2011), .CK(clk), .RN(n1507), .Q(
        \gbuff[24][16] ) );
  DFFRX1 \gbuff_reg[24][15]  ( .D(n2012), .CK(clk), .RN(n1507), .Q(
        \gbuff[24][15] ) );
  DFFRX1 \gbuff_reg[24][14]  ( .D(n2013), .CK(clk), .RN(n1507), .Q(
        \gbuff[24][14] ) );
  DFFRX1 \gbuff_reg[24][13]  ( .D(n2014), .CK(clk), .RN(n1507), .Q(
        \gbuff[24][13] ) );
  DFFRX1 \gbuff_reg[24][12]  ( .D(n2015), .CK(clk), .RN(n1507), .Q(
        \gbuff[24][12] ) );
  DFFRX1 \gbuff_reg[24][11]  ( .D(n2016), .CK(clk), .RN(n1506), .Q(
        \gbuff[24][11] ) );
  DFFRX1 \gbuff_reg[24][10]  ( .D(n2017), .CK(clk), .RN(n1506), .Q(
        \gbuff[24][10] ) );
  DFFRX1 \gbuff_reg[24][9]  ( .D(n2018), .CK(clk), .RN(n1506), .Q(
        \gbuff[24][9] ) );
  DFFRX1 \gbuff_reg[24][8]  ( .D(n2019), .CK(clk), .RN(n1506), .Q(
        \gbuff[24][8] ) );
  DFFRX1 \gbuff_reg[24][7]  ( .D(n2020), .CK(clk), .RN(n1506), .Q(
        \gbuff[24][7] ) );
  DFFRX1 \gbuff_reg[24][6]  ( .D(n2021), .CK(clk), .RN(n1506), .Q(
        \gbuff[24][6] ) );
  DFFRX1 \gbuff_reg[24][5]  ( .D(n2022), .CK(clk), .RN(n1506), .Q(
        \gbuff[24][5] ) );
  DFFRX1 \gbuff_reg[24][4]  ( .D(n2023), .CK(clk), .RN(n1506), .Q(
        \gbuff[24][4] ) );
  DFFRX1 \gbuff_reg[24][3]  ( .D(n2024), .CK(clk), .RN(n1506), .Q(
        \gbuff[24][3] ) );
  DFFRX1 \gbuff_reg[24][2]  ( .D(n2025), .CK(clk), .RN(n1506), .Q(
        \gbuff[24][2] ) );
  DFFRX1 \gbuff_reg[24][1]  ( .D(n2026), .CK(clk), .RN(n1506), .Q(
        \gbuff[24][1] ) );
  DFFRX1 \gbuff_reg[24][0]  ( .D(n2027), .CK(clk), .RN(n1506), .Q(
        \gbuff[24][0] ) );
  DFFRX1 \gbuff_reg[20][31]  ( .D(n2124), .CK(clk), .RN(n1497), .Q(
        \gbuff[20][31] ) );
  DFFRX1 \gbuff_reg[20][30]  ( .D(n2125), .CK(clk), .RN(n1497), .Q(
        \gbuff[20][30] ) );
  DFFRX1 \gbuff_reg[20][29]  ( .D(n2126), .CK(clk), .RN(n1497), .Q(
        \gbuff[20][29] ) );
  DFFRX1 \gbuff_reg[20][28]  ( .D(n2127), .CK(clk), .RN(n1497), .Q(
        \gbuff[20][28] ) );
  DFFRX1 \gbuff_reg[20][27]  ( .D(n2128), .CK(clk), .RN(n1497), .Q(
        \gbuff[20][27] ) );
  DFFRX1 \gbuff_reg[20][26]  ( .D(n2129), .CK(clk), .RN(n1497), .Q(
        \gbuff[20][26] ) );
  DFFRX1 \gbuff_reg[20][25]  ( .D(n2130), .CK(clk), .RN(n1497), .Q(
        \gbuff[20][25] ) );
  DFFRX1 \gbuff_reg[20][24]  ( .D(n2131), .CK(clk), .RN(n1497), .Q(
        \gbuff[20][24] ) );
  DFFRX1 \gbuff_reg[20][23]  ( .D(n2132), .CK(clk), .RN(n1497), .Q(
        \gbuff[20][23] ) );
  DFFRX1 \gbuff_reg[20][22]  ( .D(n2133), .CK(clk), .RN(n1497), .Q(
        \gbuff[20][22] ) );
  DFFRX1 \gbuff_reg[20][21]  ( .D(n2134), .CK(clk), .RN(n1497), .Q(
        \gbuff[20][21] ) );
  DFFRX1 \gbuff_reg[20][20]  ( .D(n2135), .CK(clk), .RN(n1497), .Q(
        \gbuff[20][20] ) );
  DFFRX1 \gbuff_reg[20][19]  ( .D(n2136), .CK(clk), .RN(n1496), .Q(
        \gbuff[20][19] ) );
  DFFRX1 \gbuff_reg[20][18]  ( .D(n2137), .CK(clk), .RN(n1496), .Q(
        \gbuff[20][18] ) );
  DFFRX1 \gbuff_reg[20][17]  ( .D(n2138), .CK(clk), .RN(n1496), .Q(
        \gbuff[20][17] ) );
  DFFRX1 \gbuff_reg[20][16]  ( .D(n2139), .CK(clk), .RN(n1496), .Q(
        \gbuff[20][16] ) );
  DFFRX1 \gbuff_reg[20][15]  ( .D(n2140), .CK(clk), .RN(n1496), .Q(
        \gbuff[20][15] ) );
  DFFRX1 \gbuff_reg[20][14]  ( .D(n2141), .CK(clk), .RN(n1496), .Q(
        \gbuff[20][14] ) );
  DFFRX1 \gbuff_reg[20][13]  ( .D(n2142), .CK(clk), .RN(n1496), .Q(
        \gbuff[20][13] ) );
  DFFRX1 \gbuff_reg[20][12]  ( .D(n2143), .CK(clk), .RN(n1496), .Q(
        \gbuff[20][12] ) );
  DFFRX1 \gbuff_reg[20][11]  ( .D(n2144), .CK(clk), .RN(n1496), .Q(
        \gbuff[20][11] ) );
  DFFRX1 \gbuff_reg[20][10]  ( .D(n2145), .CK(clk), .RN(n1496), .Q(
        \gbuff[20][10] ) );
  DFFRX1 \gbuff_reg[20][9]  ( .D(n2146), .CK(clk), .RN(n1496), .Q(
        \gbuff[20][9] ) );
  DFFRX1 \gbuff_reg[20][8]  ( .D(n2147), .CK(clk), .RN(n1496), .Q(
        \gbuff[20][8] ) );
  DFFRX1 \gbuff_reg[20][7]  ( .D(n2148), .CK(clk), .RN(n1495), .Q(
        \gbuff[20][7] ) );
  DFFRX1 \gbuff_reg[20][6]  ( .D(n2149), .CK(clk), .RN(n1495), .Q(
        \gbuff[20][6] ) );
  DFFRX1 \gbuff_reg[20][5]  ( .D(n2150), .CK(clk), .RN(n1495), .Q(
        \gbuff[20][5] ) );
  DFFRX1 \gbuff_reg[20][4]  ( .D(n2151), .CK(clk), .RN(n1495), .Q(
        \gbuff[20][4] ) );
  DFFRX1 \gbuff_reg[20][3]  ( .D(n2152), .CK(clk), .RN(n1495), .Q(
        \gbuff[20][3] ) );
  DFFRX1 \gbuff_reg[20][2]  ( .D(n2153), .CK(clk), .RN(n1495), .Q(
        \gbuff[20][2] ) );
  DFFRX1 \gbuff_reg[20][1]  ( .D(n2154), .CK(clk), .RN(n1495), .Q(
        \gbuff[20][1] ) );
  DFFRX1 \gbuff_reg[20][0]  ( .D(n2155), .CK(clk), .RN(n1495), .Q(
        \gbuff[20][0] ) );
  DFFRX1 \gbuff_reg[16][31]  ( .D(n2252), .CK(clk), .RN(n1487), .Q(
        \gbuff[16][31] ) );
  DFFRX1 \gbuff_reg[16][30]  ( .D(n2253), .CK(clk), .RN(n1487), .Q(
        \gbuff[16][30] ) );
  DFFRX1 \gbuff_reg[16][29]  ( .D(n2254), .CK(clk), .RN(n1487), .Q(
        \gbuff[16][29] ) );
  DFFRX1 \gbuff_reg[16][28]  ( .D(n2255), .CK(clk), .RN(n1487), .Q(
        \gbuff[16][28] ) );
  DFFRX1 \gbuff_reg[16][27]  ( .D(n2256), .CK(clk), .RN(n1486), .Q(
        \gbuff[16][27] ) );
  DFFRX1 \gbuff_reg[16][26]  ( .D(n2257), .CK(clk), .RN(n1486), .Q(
        \gbuff[16][26] ) );
  DFFRX1 \gbuff_reg[16][25]  ( .D(n2258), .CK(clk), .RN(n1486), .Q(
        \gbuff[16][25] ) );
  DFFRX1 \gbuff_reg[16][24]  ( .D(n2259), .CK(clk), .RN(n1486), .Q(
        \gbuff[16][24] ) );
  DFFRX1 \gbuff_reg[16][23]  ( .D(n2260), .CK(clk), .RN(n1486), .Q(
        \gbuff[16][23] ) );
  DFFRX1 \gbuff_reg[16][22]  ( .D(n2261), .CK(clk), .RN(n1486), .Q(
        \gbuff[16][22] ) );
  DFFRX1 \gbuff_reg[16][21]  ( .D(n2262), .CK(clk), .RN(n1486), .Q(
        \gbuff[16][21] ) );
  DFFRX1 \gbuff_reg[16][20]  ( .D(n2263), .CK(clk), .RN(n1486), .Q(
        \gbuff[16][20] ) );
  DFFRX1 \gbuff_reg[16][19]  ( .D(n2264), .CK(clk), .RN(n1486), .Q(
        \gbuff[16][19] ) );
  DFFRX1 \gbuff_reg[16][18]  ( .D(n2265), .CK(clk), .RN(n1486), .Q(
        \gbuff[16][18] ) );
  DFFRX1 \gbuff_reg[16][17]  ( .D(n2266), .CK(clk), .RN(n1486), .Q(
        \gbuff[16][17] ) );
  DFFRX1 \gbuff_reg[16][16]  ( .D(n2267), .CK(clk), .RN(n1486), .Q(
        \gbuff[16][16] ) );
  DFFRX1 \gbuff_reg[16][15]  ( .D(n2268), .CK(clk), .RN(n1485), .Q(
        \gbuff[16][15] ) );
  DFFRX1 \gbuff_reg[16][14]  ( .D(n2269), .CK(clk), .RN(n1485), .Q(
        \gbuff[16][14] ) );
  DFFRX1 \gbuff_reg[16][13]  ( .D(n2270), .CK(clk), .RN(n1485), .Q(
        \gbuff[16][13] ) );
  DFFRX1 \gbuff_reg[16][12]  ( .D(n2271), .CK(clk), .RN(n1485), .Q(
        \gbuff[16][12] ) );
  DFFRX1 \gbuff_reg[16][11]  ( .D(n2272), .CK(clk), .RN(n1485), .Q(
        \gbuff[16][11] ) );
  DFFRX1 \gbuff_reg[16][10]  ( .D(n2273), .CK(clk), .RN(n1485), .Q(
        \gbuff[16][10] ) );
  DFFRX1 \gbuff_reg[16][9]  ( .D(n2274), .CK(clk), .RN(n1485), .Q(
        \gbuff[16][9] ) );
  DFFRX1 \gbuff_reg[16][8]  ( .D(n2275), .CK(clk), .RN(n1485), .Q(
        \gbuff[16][8] ) );
  DFFRX1 \gbuff_reg[16][7]  ( .D(n2276), .CK(clk), .RN(n1485), .Q(
        \gbuff[16][7] ) );
  DFFRX1 \gbuff_reg[16][6]  ( .D(n2277), .CK(clk), .RN(n1485), .Q(
        \gbuff[16][6] ) );
  DFFRX1 \gbuff_reg[16][5]  ( .D(n2278), .CK(clk), .RN(n1485), .Q(
        \gbuff[16][5] ) );
  DFFRX1 \gbuff_reg[16][4]  ( .D(n2279), .CK(clk), .RN(n1485), .Q(
        \gbuff[16][4] ) );
  DFFRX1 \gbuff_reg[16][3]  ( .D(n2280), .CK(clk), .RN(n1484), .Q(
        \gbuff[16][3] ) );
  DFFRX1 \gbuff_reg[16][2]  ( .D(n2281), .CK(clk), .RN(n1484), .Q(
        \gbuff[16][2] ) );
  DFFRX1 \gbuff_reg[16][1]  ( .D(n2282), .CK(clk), .RN(n1484), .Q(
        \gbuff[16][1] ) );
  DFFRX1 \gbuff_reg[16][0]  ( .D(n2283), .CK(clk), .RN(n1484), .Q(
        \gbuff[16][0] ) );
  DFFRX1 \gbuff_reg[12][31]  ( .D(n2380), .CK(clk), .RN(n1476), .Q(
        \gbuff[12][31] ) );
  DFFRX1 \gbuff_reg[12][30]  ( .D(n2381), .CK(clk), .RN(n1476), .Q(
        \gbuff[12][30] ) );
  DFFRX1 \gbuff_reg[12][29]  ( .D(n2382), .CK(clk), .RN(n1476), .Q(
        \gbuff[12][29] ) );
  DFFRX1 \gbuff_reg[12][28]  ( .D(n2383), .CK(clk), .RN(n1476), .Q(
        \gbuff[12][28] ) );
  DFFRX1 \gbuff_reg[12][27]  ( .D(n2384), .CK(clk), .RN(n1476), .Q(
        \gbuff[12][27] ) );
  DFFRX1 \gbuff_reg[12][26]  ( .D(n2385), .CK(clk), .RN(n1476), .Q(
        \gbuff[12][26] ) );
  DFFRX1 \gbuff_reg[12][25]  ( .D(n2386), .CK(clk), .RN(n1476), .Q(
        \gbuff[12][25] ) );
  DFFRX1 \gbuff_reg[12][24]  ( .D(n2387), .CK(clk), .RN(n1476), .Q(
        \gbuff[12][24] ) );
  DFFRX1 \gbuff_reg[12][23]  ( .D(n2388), .CK(clk), .RN(n1475), .Q(
        \gbuff[12][23] ) );
  DFFRX1 \gbuff_reg[12][22]  ( .D(n2389), .CK(clk), .RN(n1475), .Q(
        \gbuff[12][22] ) );
  DFFRX1 \gbuff_reg[12][21]  ( .D(n2390), .CK(clk), .RN(n1475), .Q(
        \gbuff[12][21] ) );
  DFFRX1 \gbuff_reg[12][20]  ( .D(n2391), .CK(clk), .RN(n1475), .Q(
        \gbuff[12][20] ) );
  DFFRX1 \gbuff_reg[12][19]  ( .D(n2392), .CK(clk), .RN(n1475), .Q(
        \gbuff[12][19] ) );
  DFFRX1 \gbuff_reg[12][18]  ( .D(n2393), .CK(clk), .RN(n1475), .Q(
        \gbuff[12][18] ) );
  DFFRX1 \gbuff_reg[12][17]  ( .D(n2394), .CK(clk), .RN(n1475), .Q(
        \gbuff[12][17] ) );
  DFFRX1 \gbuff_reg[12][16]  ( .D(n2395), .CK(clk), .RN(n1475), .Q(
        \gbuff[12][16] ) );
  DFFRX1 \gbuff_reg[12][15]  ( .D(n2396), .CK(clk), .RN(n1475), .Q(
        \gbuff[12][15] ) );
  DFFRX1 \gbuff_reg[12][14]  ( .D(n2397), .CK(clk), .RN(n1475), .Q(
        \gbuff[12][14] ) );
  DFFRX1 \gbuff_reg[12][13]  ( .D(n2398), .CK(clk), .RN(n1475), .Q(
        \gbuff[12][13] ) );
  DFFRX1 \gbuff_reg[12][12]  ( .D(n2399), .CK(clk), .RN(n1475), .Q(
        \gbuff[12][12] ) );
  DFFRX1 \gbuff_reg[12][11]  ( .D(n2400), .CK(clk), .RN(n1474), .Q(
        \gbuff[12][11] ) );
  DFFRX1 \gbuff_reg[12][10]  ( .D(n2401), .CK(clk), .RN(n1474), .Q(
        \gbuff[12][10] ) );
  DFFRX1 \gbuff_reg[12][9]  ( .D(n2402), .CK(clk), .RN(n1474), .Q(
        \gbuff[12][9] ) );
  DFFRX1 \gbuff_reg[12][8]  ( .D(n2403), .CK(clk), .RN(n1474), .Q(
        \gbuff[12][8] ) );
  DFFRX1 \gbuff_reg[12][7]  ( .D(n2404), .CK(clk), .RN(n1474), .Q(
        \gbuff[12][7] ) );
  DFFRX1 \gbuff_reg[12][6]  ( .D(n2405), .CK(clk), .RN(n1474), .Q(
        \gbuff[12][6] ) );
  DFFRX1 \gbuff_reg[12][5]  ( .D(n2406), .CK(clk), .RN(n1474), .Q(
        \gbuff[12][5] ) );
  DFFRX1 \gbuff_reg[12][4]  ( .D(n2407), .CK(clk), .RN(n1474), .Q(
        \gbuff[12][4] ) );
  DFFRX1 \gbuff_reg[12][3]  ( .D(n2408), .CK(clk), .RN(n1474), .Q(
        \gbuff[12][3] ) );
  DFFRX1 \gbuff_reg[12][2]  ( .D(n2409), .CK(clk), .RN(n1474), .Q(
        \gbuff[12][2] ) );
  DFFRX1 \gbuff_reg[12][1]  ( .D(n2410), .CK(clk), .RN(n1474), .Q(
        \gbuff[12][1] ) );
  DFFRX1 \gbuff_reg[12][0]  ( .D(n2411), .CK(clk), .RN(n1474), .Q(
        \gbuff[12][0] ) );
  DFFRX1 \gbuff_reg[8][31]  ( .D(n2508), .CK(clk), .RN(n1465), .Q(
        \gbuff[8][31] ) );
  DFFRX1 \gbuff_reg[8][30]  ( .D(n2509), .CK(clk), .RN(n1465), .Q(
        \gbuff[8][30] ) );
  DFFRX1 \gbuff_reg[8][29]  ( .D(n2510), .CK(clk), .RN(n1465), .Q(
        \gbuff[8][29] ) );
  DFFRX1 \gbuff_reg[8][28]  ( .D(n2511), .CK(clk), .RN(n1465), .Q(
        \gbuff[8][28] ) );
  DFFRX1 \gbuff_reg[8][27]  ( .D(n2512), .CK(clk), .RN(n1465), .Q(
        \gbuff[8][27] ) );
  DFFRX1 \gbuff_reg[8][26]  ( .D(n2513), .CK(clk), .RN(n1465), .Q(
        \gbuff[8][26] ) );
  DFFRX1 \gbuff_reg[8][25]  ( .D(n2514), .CK(clk), .RN(n1465), .Q(
        \gbuff[8][25] ) );
  DFFRX1 \gbuff_reg[8][24]  ( .D(n2515), .CK(clk), .RN(n1465), .Q(
        \gbuff[8][24] ) );
  DFFRX1 \gbuff_reg[8][23]  ( .D(n2516), .CK(clk), .RN(n1465), .Q(
        \gbuff[8][23] ) );
  DFFRX1 \gbuff_reg[8][22]  ( .D(n2517), .CK(clk), .RN(n1465), .Q(
        \gbuff[8][22] ) );
  DFFRX1 \gbuff_reg[8][21]  ( .D(n2518), .CK(clk), .RN(n1465), .Q(
        \gbuff[8][21] ) );
  DFFRX1 \gbuff_reg[8][20]  ( .D(n2519), .CK(clk), .RN(n1465), .Q(
        \gbuff[8][20] ) );
  DFFRX1 \gbuff_reg[8][19]  ( .D(n2520), .CK(clk), .RN(n1464), .Q(
        \gbuff[8][19] ) );
  DFFRX1 \gbuff_reg[8][18]  ( .D(n2521), .CK(clk), .RN(n1464), .Q(
        \gbuff[8][18] ) );
  DFFRX1 \gbuff_reg[8][17]  ( .D(n2522), .CK(clk), .RN(n1464), .Q(
        \gbuff[8][17] ) );
  DFFRX1 \gbuff_reg[8][16]  ( .D(n2523), .CK(clk), .RN(n1464), .Q(
        \gbuff[8][16] ) );
  DFFRX1 \gbuff_reg[8][15]  ( .D(n2524), .CK(clk), .RN(n1464), .Q(
        \gbuff[8][15] ) );
  DFFRX1 \gbuff_reg[8][14]  ( .D(n2525), .CK(clk), .RN(n1464), .Q(
        \gbuff[8][14] ) );
  DFFRX1 \gbuff_reg[8][13]  ( .D(n2526), .CK(clk), .RN(n1464), .Q(
        \gbuff[8][13] ) );
  DFFRX1 \gbuff_reg[8][12]  ( .D(n2527), .CK(clk), .RN(n1464), .Q(
        \gbuff[8][12] ) );
  DFFRX1 \gbuff_reg[8][11]  ( .D(n2528), .CK(clk), .RN(n1464), .Q(
        \gbuff[8][11] ) );
  DFFRX1 \gbuff_reg[8][10]  ( .D(n2529), .CK(clk), .RN(n1464), .Q(
        \gbuff[8][10] ) );
  DFFRX1 \gbuff_reg[8][9]  ( .D(n2530), .CK(clk), .RN(n1464), .Q(\gbuff[8][9] ) );
  DFFRX1 \gbuff_reg[8][8]  ( .D(n2531), .CK(clk), .RN(n1464), .Q(\gbuff[8][8] ) );
  DFFRX1 \gbuff_reg[8][7]  ( .D(n2532), .CK(clk), .RN(n1463), .Q(\gbuff[8][7] ) );
  DFFRX1 \gbuff_reg[8][6]  ( .D(n2533), .CK(clk), .RN(n1463), .Q(\gbuff[8][6] ) );
  DFFRX1 \gbuff_reg[8][5]  ( .D(n2534), .CK(clk), .RN(n1463), .Q(\gbuff[8][5] ) );
  DFFRX1 \gbuff_reg[8][4]  ( .D(n2535), .CK(clk), .RN(n1463), .Q(\gbuff[8][4] ) );
  DFFRX1 \gbuff_reg[8][3]  ( .D(n2536), .CK(clk), .RN(n1463), .Q(\gbuff[8][3] ) );
  DFFRX1 \gbuff_reg[8][2]  ( .D(n2537), .CK(clk), .RN(n1463), .Q(\gbuff[8][2] ) );
  DFFRX1 \gbuff_reg[8][1]  ( .D(n2538), .CK(clk), .RN(n1463), .Q(\gbuff[8][1] ) );
  DFFRX1 \gbuff_reg[8][0]  ( .D(n2539), .CK(clk), .RN(n1463), .Q(\gbuff[8][0] ) );
  DFFRX1 \gbuff_reg[4][31]  ( .D(n2636), .CK(clk), .RN(n1455), .Q(
        \gbuff[4][31] ) );
  DFFRX1 \gbuff_reg[4][30]  ( .D(n2637), .CK(clk), .RN(n1455), .Q(
        \gbuff[4][30] ) );
  DFFRX1 \gbuff_reg[4][29]  ( .D(n2638), .CK(clk), .RN(n1455), .Q(
        \gbuff[4][29] ) );
  DFFRX1 \gbuff_reg[4][28]  ( .D(n2639), .CK(clk), .RN(n1455), .Q(
        \gbuff[4][28] ) );
  DFFRX1 \gbuff_reg[4][27]  ( .D(n2640), .CK(clk), .RN(n1454), .Q(
        \gbuff[4][27] ) );
  DFFRX1 \gbuff_reg[4][26]  ( .D(n2641), .CK(clk), .RN(n1454), .Q(
        \gbuff[4][26] ) );
  DFFRX1 \gbuff_reg[4][25]  ( .D(n2642), .CK(clk), .RN(n1454), .Q(
        \gbuff[4][25] ) );
  DFFRX1 \gbuff_reg[4][24]  ( .D(n2643), .CK(clk), .RN(n1454), .Q(
        \gbuff[4][24] ) );
  DFFRX1 \gbuff_reg[4][23]  ( .D(n2644), .CK(clk), .RN(n1454), .Q(
        \gbuff[4][23] ) );
  DFFRX1 \gbuff_reg[4][22]  ( .D(n2645), .CK(clk), .RN(n1454), .Q(
        \gbuff[4][22] ) );
  DFFRX1 \gbuff_reg[4][21]  ( .D(n2646), .CK(clk), .RN(n1454), .Q(
        \gbuff[4][21] ) );
  DFFRX1 \gbuff_reg[4][20]  ( .D(n2647), .CK(clk), .RN(n1454), .Q(
        \gbuff[4][20] ) );
  DFFRX1 \gbuff_reg[4][19]  ( .D(n2648), .CK(clk), .RN(n1454), .Q(
        \gbuff[4][19] ) );
  DFFRX1 \gbuff_reg[4][18]  ( .D(n2649), .CK(clk), .RN(n1454), .Q(
        \gbuff[4][18] ) );
  DFFRX1 \gbuff_reg[4][17]  ( .D(n2650), .CK(clk), .RN(n1454), .Q(
        \gbuff[4][17] ) );
  DFFRX1 \gbuff_reg[4][16]  ( .D(n2651), .CK(clk), .RN(n1454), .Q(
        \gbuff[4][16] ) );
  DFFRX1 \gbuff_reg[4][15]  ( .D(n2652), .CK(clk), .RN(n1453), .Q(
        \gbuff[4][15] ) );
  DFFRX1 \gbuff_reg[4][14]  ( .D(n2653), .CK(clk), .RN(n1453), .Q(
        \gbuff[4][14] ) );
  DFFRX1 \gbuff_reg[4][13]  ( .D(n2654), .CK(clk), .RN(n1453), .Q(
        \gbuff[4][13] ) );
  DFFRX1 \gbuff_reg[4][12]  ( .D(n2655), .CK(clk), .RN(n1453), .Q(
        \gbuff[4][12] ) );
  DFFRX1 \gbuff_reg[4][11]  ( .D(n2656), .CK(clk), .RN(n1453), .Q(
        \gbuff[4][11] ) );
  DFFRX1 \gbuff_reg[4][10]  ( .D(n2657), .CK(clk), .RN(n1453), .Q(
        \gbuff[4][10] ) );
  DFFRX1 \gbuff_reg[4][9]  ( .D(n2658), .CK(clk), .RN(n1453), .Q(\gbuff[4][9] ) );
  DFFRX1 \gbuff_reg[4][8]  ( .D(n2659), .CK(clk), .RN(n1453), .Q(\gbuff[4][8] ) );
  DFFRX1 \gbuff_reg[4][7]  ( .D(n2660), .CK(clk), .RN(n1453), .Q(\gbuff[4][7] ) );
  DFFRX1 \gbuff_reg[4][6]  ( .D(n2661), .CK(clk), .RN(n1453), .Q(\gbuff[4][6] ) );
  DFFRX1 \gbuff_reg[4][5]  ( .D(n2662), .CK(clk), .RN(n1453), .Q(\gbuff[4][5] ) );
  DFFRX1 \gbuff_reg[4][4]  ( .D(n2663), .CK(clk), .RN(n1453), .Q(\gbuff[4][4] ) );
  DFFRX1 \gbuff_reg[4][3]  ( .D(n2664), .CK(clk), .RN(n1452), .Q(\gbuff[4][3] ) );
  DFFRX1 \gbuff_reg[4][2]  ( .D(n2665), .CK(clk), .RN(n1452), .Q(\gbuff[4][2] ) );
  DFFRX1 \gbuff_reg[4][1]  ( .D(n2666), .CK(clk), .RN(n1452), .Q(\gbuff[4][1] ) );
  DFFRX1 \gbuff_reg[4][0]  ( .D(n2667), .CK(clk), .RN(n1452), .Q(\gbuff[4][0] ) );
  DFFRX1 \gbuff_reg[0][31]  ( .D(n2764), .CK(clk), .RN(n1444), .Q(
        \gbuff[0][31] ) );
  DFFRX1 \gbuff_reg[0][30]  ( .D(n2765), .CK(clk), .RN(n1444), .Q(
        \gbuff[0][30] ) );
  DFFRX1 \gbuff_reg[0][29]  ( .D(n2766), .CK(clk), .RN(n1444), .Q(
        \gbuff[0][29] ) );
  DFFRX1 \gbuff_reg[0][28]  ( .D(n2767), .CK(clk), .RN(n1444), .Q(
        \gbuff[0][28] ) );
  DFFRX1 \gbuff_reg[0][27]  ( .D(n2768), .CK(clk), .RN(n1444), .Q(
        \gbuff[0][27] ) );
  DFFRX1 \gbuff_reg[0][26]  ( .D(n2769), .CK(clk), .RN(n1444), .Q(
        \gbuff[0][26] ) );
  DFFRX1 \gbuff_reg[0][25]  ( .D(n2770), .CK(clk), .RN(n1444), .Q(
        \gbuff[0][25] ) );
  DFFRX1 \gbuff_reg[0][24]  ( .D(n2771), .CK(clk), .RN(n1444), .Q(
        \gbuff[0][24] ) );
  DFFRX1 \gbuff_reg[0][23]  ( .D(n2772), .CK(clk), .RN(n1443), .Q(
        \gbuff[0][23] ) );
  DFFRX1 \gbuff_reg[0][22]  ( .D(n2773), .CK(clk), .RN(n1443), .Q(
        \gbuff[0][22] ) );
  DFFRX1 \gbuff_reg[0][21]  ( .D(n2774), .CK(clk), .RN(n1443), .Q(
        \gbuff[0][21] ) );
  DFFRX1 \gbuff_reg[0][20]  ( .D(n2775), .CK(clk), .RN(n1443), .Q(
        \gbuff[0][20] ) );
  DFFRX1 \gbuff_reg[0][19]  ( .D(n2776), .CK(clk), .RN(n1443), .Q(
        \gbuff[0][19] ) );
  DFFRX1 \gbuff_reg[0][18]  ( .D(n2777), .CK(clk), .RN(n1443), .Q(
        \gbuff[0][18] ) );
  DFFRX1 \gbuff_reg[0][17]  ( .D(n2778), .CK(clk), .RN(n1443), .Q(
        \gbuff[0][17] ) );
  DFFRX1 \gbuff_reg[0][16]  ( .D(n2779), .CK(clk), .RN(n1443), .Q(
        \gbuff[0][16] ) );
  DFFRX1 \gbuff_reg[0][15]  ( .D(n2780), .CK(clk), .RN(n1443), .Q(
        \gbuff[0][15] ) );
  DFFRX1 \gbuff_reg[0][14]  ( .D(n2781), .CK(clk), .RN(n1443), .Q(
        \gbuff[0][14] ) );
  DFFRX1 \gbuff_reg[0][13]  ( .D(n2782), .CK(clk), .RN(n1443), .Q(
        \gbuff[0][13] ) );
  DFFRX1 \gbuff_reg[0][12]  ( .D(n2783), .CK(clk), .RN(n1443), .Q(
        \gbuff[0][12] ) );
  DFFRX1 \gbuff_reg[0][11]  ( .D(n2784), .CK(clk), .RN(n1442), .Q(
        \gbuff[0][11] ) );
  DFFRX1 \gbuff_reg[0][10]  ( .D(n2785), .CK(clk), .RN(n1442), .Q(
        \gbuff[0][10] ) );
  DFFRX1 \gbuff_reg[0][9]  ( .D(n2786), .CK(clk), .RN(n1442), .Q(\gbuff[0][9] ) );
  DFFRX1 \gbuff_reg[0][8]  ( .D(n2787), .CK(clk), .RN(n1442), .Q(\gbuff[0][8] ) );
  DFFRX1 \gbuff_reg[0][7]  ( .D(n2788), .CK(clk), .RN(n1442), .Q(\gbuff[0][7] ) );
  DFFRX1 \gbuff_reg[0][6]  ( .D(n2789), .CK(clk), .RN(n1442), .Q(\gbuff[0][6] ) );
  DFFRX1 \gbuff_reg[0][5]  ( .D(n2790), .CK(clk), .RN(n1442), .Q(\gbuff[0][5] ) );
  DFFRX1 \gbuff_reg[0][4]  ( .D(n2791), .CK(clk), .RN(n1442), .Q(\gbuff[0][4] ) );
  DFFRX1 \gbuff_reg[0][3]  ( .D(n2792), .CK(clk), .RN(n1442), .Q(\gbuff[0][3] ) );
  DFFRX1 \gbuff_reg[0][2]  ( .D(n2793), .CK(clk), .RN(n1442), .Q(\gbuff[0][2] ) );
  DFFRX1 \gbuff_reg[0][1]  ( .D(n2794), .CK(clk), .RN(n1442), .Q(\gbuff[0][1] ) );
  DFFRX1 \gbuff_reg[0][0]  ( .D(n2795), .CK(clk), .RN(n1442), .Q(\gbuff[0][0] ) );
  DFFRX1 \gbuff_reg[30][31]  ( .D(n1804), .CK(clk), .RN(n1524), .Q(
        \gbuff[30][31] ) );
  DFFRX1 \gbuff_reg[30][30]  ( .D(n1805), .CK(clk), .RN(n1524), .Q(
        \gbuff[30][30] ) );
  DFFRX1 \gbuff_reg[30][29]  ( .D(n1806), .CK(clk), .RN(n1524), .Q(
        \gbuff[30][29] ) );
  DFFRX1 \gbuff_reg[30][28]  ( .D(n1807), .CK(clk), .RN(n1524), .Q(
        \gbuff[30][28] ) );
  DFFRX1 \gbuff_reg[30][27]  ( .D(n1808), .CK(clk), .RN(n1524), .Q(
        \gbuff[30][27] ) );
  DFFRX1 \gbuff_reg[30][26]  ( .D(n1809), .CK(clk), .RN(n1524), .Q(
        \gbuff[30][26] ) );
  DFFRX1 \gbuff_reg[30][25]  ( .D(n1810), .CK(clk), .RN(n1524), .Q(
        \gbuff[30][25] ) );
  DFFRX1 \gbuff_reg[30][24]  ( .D(n1811), .CK(clk), .RN(n1524), .Q(
        \gbuff[30][24] ) );
  DFFRX1 \gbuff_reg[30][23]  ( .D(n1812), .CK(clk), .RN(n1523), .Q(
        \gbuff[30][23] ) );
  DFFRX1 \gbuff_reg[30][22]  ( .D(n1813), .CK(clk), .RN(n1523), .Q(
        \gbuff[30][22] ) );
  DFFRX1 \gbuff_reg[30][21]  ( .D(n1814), .CK(clk), .RN(n1523), .Q(
        \gbuff[30][21] ) );
  DFFRX1 \gbuff_reg[30][20]  ( .D(n1815), .CK(clk), .RN(n1523), .Q(
        \gbuff[30][20] ) );
  DFFRX1 \gbuff_reg[30][19]  ( .D(n1816), .CK(clk), .RN(n1523), .Q(
        \gbuff[30][19] ) );
  DFFRX1 \gbuff_reg[30][18]  ( .D(n1817), .CK(clk), .RN(n1523), .Q(
        \gbuff[30][18] ) );
  DFFRX1 \gbuff_reg[30][17]  ( .D(n1818), .CK(clk), .RN(n1523), .Q(
        \gbuff[30][17] ) );
  DFFRX1 \gbuff_reg[30][16]  ( .D(n1819), .CK(clk), .RN(n1523), .Q(
        \gbuff[30][16] ) );
  DFFRX1 \gbuff_reg[30][15]  ( .D(n1820), .CK(clk), .RN(n1523), .Q(
        \gbuff[30][15] ) );
  DFFRX1 \gbuff_reg[30][14]  ( .D(n1821), .CK(clk), .RN(n1523), .Q(
        \gbuff[30][14] ) );
  DFFRX1 \gbuff_reg[30][13]  ( .D(n1822), .CK(clk), .RN(n1523), .Q(
        \gbuff[30][13] ) );
  DFFRX1 \gbuff_reg[30][12]  ( .D(n1823), .CK(clk), .RN(n1523), .Q(
        \gbuff[30][12] ) );
  DFFRX1 \gbuff_reg[30][11]  ( .D(n1824), .CK(clk), .RN(n1522), .Q(
        \gbuff[30][11] ) );
  DFFRX1 \gbuff_reg[30][10]  ( .D(n1825), .CK(clk), .RN(n1522), .Q(
        \gbuff[30][10] ) );
  DFFRX1 \gbuff_reg[30][9]  ( .D(n1826), .CK(clk), .RN(n1522), .Q(
        \gbuff[30][9] ) );
  DFFRX1 \gbuff_reg[30][8]  ( .D(n1827), .CK(clk), .RN(n1522), .Q(
        \gbuff[30][8] ) );
  DFFRX1 \gbuff_reg[30][7]  ( .D(n1828), .CK(clk), .RN(n1522), .Q(
        \gbuff[30][7] ) );
  DFFRX1 \gbuff_reg[30][6]  ( .D(n1829), .CK(clk), .RN(n1522), .Q(
        \gbuff[30][6] ) );
  DFFRX1 \gbuff_reg[30][5]  ( .D(n1830), .CK(clk), .RN(n1522), .Q(
        \gbuff[30][5] ) );
  DFFRX1 \gbuff_reg[30][4]  ( .D(n1831), .CK(clk), .RN(n1522), .Q(
        \gbuff[30][4] ) );
  DFFRX1 \gbuff_reg[30][3]  ( .D(n1832), .CK(clk), .RN(n1522), .Q(
        \gbuff[30][3] ) );
  DFFRX1 \gbuff_reg[30][2]  ( .D(n1833), .CK(clk), .RN(n1522), .Q(
        \gbuff[30][2] ) );
  DFFRX1 \gbuff_reg[30][1]  ( .D(n1834), .CK(clk), .RN(n1522), .Q(
        \gbuff[30][1] ) );
  DFFRX1 \gbuff_reg[30][0]  ( .D(n1835), .CK(clk), .RN(n1522), .Q(
        \gbuff[30][0] ) );
  DFFRX1 \gbuff_reg[26][31]  ( .D(n1932), .CK(clk), .RN(n1513), .Q(
        \gbuff[26][31] ) );
  DFFRX1 \gbuff_reg[26][30]  ( .D(n1933), .CK(clk), .RN(n1513), .Q(
        \gbuff[26][30] ) );
  DFFRX1 \gbuff_reg[26][29]  ( .D(n1934), .CK(clk), .RN(n1513), .Q(
        \gbuff[26][29] ) );
  DFFRX1 \gbuff_reg[26][28]  ( .D(n1935), .CK(clk), .RN(n1513), .Q(
        \gbuff[26][28] ) );
  DFFRX1 \gbuff_reg[26][27]  ( .D(n1936), .CK(clk), .RN(n1513), .Q(
        \gbuff[26][27] ) );
  DFFRX1 \gbuff_reg[26][26]  ( .D(n1937), .CK(clk), .RN(n1513), .Q(
        \gbuff[26][26] ) );
  DFFRX1 \gbuff_reg[26][25]  ( .D(n1938), .CK(clk), .RN(n1513), .Q(
        \gbuff[26][25] ) );
  DFFRX1 \gbuff_reg[26][24]  ( .D(n1939), .CK(clk), .RN(n1513), .Q(
        \gbuff[26][24] ) );
  DFFRX1 \gbuff_reg[26][23]  ( .D(n1940), .CK(clk), .RN(n1513), .Q(
        \gbuff[26][23] ) );
  DFFRX1 \gbuff_reg[26][22]  ( .D(n1941), .CK(clk), .RN(n1513), .Q(
        \gbuff[26][22] ) );
  DFFRX1 \gbuff_reg[26][21]  ( .D(n1942), .CK(clk), .RN(n1513), .Q(
        \gbuff[26][21] ) );
  DFFRX1 \gbuff_reg[26][20]  ( .D(n1943), .CK(clk), .RN(n1513), .Q(
        \gbuff[26][20] ) );
  DFFRX1 \gbuff_reg[26][19]  ( .D(n1944), .CK(clk), .RN(n1512), .Q(
        \gbuff[26][19] ) );
  DFFRX1 \gbuff_reg[26][18]  ( .D(n1945), .CK(clk), .RN(n1512), .Q(
        \gbuff[26][18] ) );
  DFFRX1 \gbuff_reg[26][17]  ( .D(n1946), .CK(clk), .RN(n1512), .Q(
        \gbuff[26][17] ) );
  DFFRX1 \gbuff_reg[26][16]  ( .D(n1947), .CK(clk), .RN(n1512), .Q(
        \gbuff[26][16] ) );
  DFFRX1 \gbuff_reg[26][15]  ( .D(n1948), .CK(clk), .RN(n1512), .Q(
        \gbuff[26][15] ) );
  DFFRX1 \gbuff_reg[26][14]  ( .D(n1949), .CK(clk), .RN(n1512), .Q(
        \gbuff[26][14] ) );
  DFFRX1 \gbuff_reg[26][13]  ( .D(n1950), .CK(clk), .RN(n1512), .Q(
        \gbuff[26][13] ) );
  DFFRX1 \gbuff_reg[26][12]  ( .D(n1951), .CK(clk), .RN(n1512), .Q(
        \gbuff[26][12] ) );
  DFFRX1 \gbuff_reg[26][11]  ( .D(n1952), .CK(clk), .RN(n1512), .Q(
        \gbuff[26][11] ) );
  DFFRX1 \gbuff_reg[26][10]  ( .D(n1953), .CK(clk), .RN(n1512), .Q(
        \gbuff[26][10] ) );
  DFFRX1 \gbuff_reg[26][9]  ( .D(n1954), .CK(clk), .RN(n1512), .Q(
        \gbuff[26][9] ) );
  DFFRX1 \gbuff_reg[26][8]  ( .D(n1955), .CK(clk), .RN(n1512), .Q(
        \gbuff[26][8] ) );
  DFFRX1 \gbuff_reg[26][7]  ( .D(n1956), .CK(clk), .RN(n1511), .Q(
        \gbuff[26][7] ) );
  DFFRX1 \gbuff_reg[26][6]  ( .D(n1957), .CK(clk), .RN(n1511), .Q(
        \gbuff[26][6] ) );
  DFFRX1 \gbuff_reg[26][5]  ( .D(n1958), .CK(clk), .RN(n1511), .Q(
        \gbuff[26][5] ) );
  DFFRX1 \gbuff_reg[26][4]  ( .D(n1959), .CK(clk), .RN(n1511), .Q(
        \gbuff[26][4] ) );
  DFFRX1 \gbuff_reg[26][3]  ( .D(n1960), .CK(clk), .RN(n1511), .Q(
        \gbuff[26][3] ) );
  DFFRX1 \gbuff_reg[26][2]  ( .D(n1961), .CK(clk), .RN(n1511), .Q(
        \gbuff[26][2] ) );
  DFFRX1 \gbuff_reg[26][1]  ( .D(n1962), .CK(clk), .RN(n1511), .Q(
        \gbuff[26][1] ) );
  DFFRX1 \gbuff_reg[26][0]  ( .D(n1963), .CK(clk), .RN(n1511), .Q(
        \gbuff[26][0] ) );
  DFFRX1 \gbuff_reg[22][31]  ( .D(n2060), .CK(clk), .RN(n1503), .Q(
        \gbuff[22][31] ) );
  DFFRX1 \gbuff_reg[22][30]  ( .D(n2061), .CK(clk), .RN(n1503), .Q(
        \gbuff[22][30] ) );
  DFFRX1 \gbuff_reg[22][29]  ( .D(n2062), .CK(clk), .RN(n1503), .Q(
        \gbuff[22][29] ) );
  DFFRX1 \gbuff_reg[22][28]  ( .D(n2063), .CK(clk), .RN(n1503), .Q(
        \gbuff[22][28] ) );
  DFFRX1 \gbuff_reg[22][27]  ( .D(n2064), .CK(clk), .RN(n1502), .Q(
        \gbuff[22][27] ) );
  DFFRX1 \gbuff_reg[22][26]  ( .D(n2065), .CK(clk), .RN(n1502), .Q(
        \gbuff[22][26] ) );
  DFFRX1 \gbuff_reg[22][25]  ( .D(n2066), .CK(clk), .RN(n1502), .Q(
        \gbuff[22][25] ) );
  DFFRX1 \gbuff_reg[22][24]  ( .D(n2067), .CK(clk), .RN(n1502), .Q(
        \gbuff[22][24] ) );
  DFFRX1 \gbuff_reg[22][23]  ( .D(n2068), .CK(clk), .RN(n1502), .Q(
        \gbuff[22][23] ) );
  DFFRX1 \gbuff_reg[22][22]  ( .D(n2069), .CK(clk), .RN(n1502), .Q(
        \gbuff[22][22] ) );
  DFFRX1 \gbuff_reg[22][21]  ( .D(n2070), .CK(clk), .RN(n1502), .Q(
        \gbuff[22][21] ) );
  DFFRX1 \gbuff_reg[22][20]  ( .D(n2071), .CK(clk), .RN(n1502), .Q(
        \gbuff[22][20] ) );
  DFFRX1 \gbuff_reg[22][19]  ( .D(n2072), .CK(clk), .RN(n1502), .Q(
        \gbuff[22][19] ) );
  DFFRX1 \gbuff_reg[22][18]  ( .D(n2073), .CK(clk), .RN(n1502), .Q(
        \gbuff[22][18] ) );
  DFFRX1 \gbuff_reg[22][17]  ( .D(n2074), .CK(clk), .RN(n1502), .Q(
        \gbuff[22][17] ) );
  DFFRX1 \gbuff_reg[22][16]  ( .D(n2075), .CK(clk), .RN(n1502), .Q(
        \gbuff[22][16] ) );
  DFFRX1 \gbuff_reg[22][15]  ( .D(n2076), .CK(clk), .RN(n1501), .Q(
        \gbuff[22][15] ) );
  DFFRX1 \gbuff_reg[22][14]  ( .D(n2077), .CK(clk), .RN(n1501), .Q(
        \gbuff[22][14] ) );
  DFFRX1 \gbuff_reg[22][13]  ( .D(n2078), .CK(clk), .RN(n1501), .Q(
        \gbuff[22][13] ) );
  DFFRX1 \gbuff_reg[22][12]  ( .D(n2079), .CK(clk), .RN(n1501), .Q(
        \gbuff[22][12] ) );
  DFFRX1 \gbuff_reg[22][11]  ( .D(n2080), .CK(clk), .RN(n1501), .Q(
        \gbuff[22][11] ) );
  DFFRX1 \gbuff_reg[22][10]  ( .D(n2081), .CK(clk), .RN(n1501), .Q(
        \gbuff[22][10] ) );
  DFFRX1 \gbuff_reg[22][9]  ( .D(n2082), .CK(clk), .RN(n1501), .Q(
        \gbuff[22][9] ) );
  DFFRX1 \gbuff_reg[22][8]  ( .D(n2083), .CK(clk), .RN(n1501), .Q(
        \gbuff[22][8] ) );
  DFFRX1 \gbuff_reg[22][7]  ( .D(n2084), .CK(clk), .RN(n1501), .Q(
        \gbuff[22][7] ) );
  DFFRX1 \gbuff_reg[22][6]  ( .D(n2085), .CK(clk), .RN(n1501), .Q(
        \gbuff[22][6] ) );
  DFFRX1 \gbuff_reg[22][5]  ( .D(n2086), .CK(clk), .RN(n1501), .Q(
        \gbuff[22][5] ) );
  DFFRX1 \gbuff_reg[22][4]  ( .D(n2087), .CK(clk), .RN(n1501), .Q(
        \gbuff[22][4] ) );
  DFFRX1 \gbuff_reg[22][3]  ( .D(n2088), .CK(clk), .RN(n1500), .Q(
        \gbuff[22][3] ) );
  DFFRX1 \gbuff_reg[22][2]  ( .D(n2089), .CK(clk), .RN(n1500), .Q(
        \gbuff[22][2] ) );
  DFFRX1 \gbuff_reg[22][1]  ( .D(n2090), .CK(clk), .RN(n1500), .Q(
        \gbuff[22][1] ) );
  DFFRX1 \gbuff_reg[22][0]  ( .D(n2091), .CK(clk), .RN(n1500), .Q(
        \gbuff[22][0] ) );
  DFFRX1 \gbuff_reg[18][31]  ( .D(n2188), .CK(clk), .RN(n1492), .Q(
        \gbuff[18][31] ) );
  DFFRX1 \gbuff_reg[18][30]  ( .D(n2189), .CK(clk), .RN(n1492), .Q(
        \gbuff[18][30] ) );
  DFFRX1 \gbuff_reg[18][29]  ( .D(n2190), .CK(clk), .RN(n1492), .Q(
        \gbuff[18][29] ) );
  DFFRX1 \gbuff_reg[18][28]  ( .D(n2191), .CK(clk), .RN(n1492), .Q(
        \gbuff[18][28] ) );
  DFFRX1 \gbuff_reg[18][27]  ( .D(n2192), .CK(clk), .RN(n1492), .Q(
        \gbuff[18][27] ) );
  DFFRX1 \gbuff_reg[18][26]  ( .D(n2193), .CK(clk), .RN(n1492), .Q(
        \gbuff[18][26] ) );
  DFFRX1 \gbuff_reg[18][25]  ( .D(n2194), .CK(clk), .RN(n1492), .Q(
        \gbuff[18][25] ) );
  DFFRX1 \gbuff_reg[18][24]  ( .D(n2195), .CK(clk), .RN(n1492), .Q(
        \gbuff[18][24] ) );
  DFFRX1 \gbuff_reg[18][23]  ( .D(n2196), .CK(clk), .RN(n1491), .Q(
        \gbuff[18][23] ) );
  DFFRX1 \gbuff_reg[18][22]  ( .D(n2197), .CK(clk), .RN(n1491), .Q(
        \gbuff[18][22] ) );
  DFFRX1 \gbuff_reg[18][21]  ( .D(n2198), .CK(clk), .RN(n1491), .Q(
        \gbuff[18][21] ) );
  DFFRX1 \gbuff_reg[18][20]  ( .D(n2199), .CK(clk), .RN(n1491), .Q(
        \gbuff[18][20] ) );
  DFFRX1 \gbuff_reg[18][19]  ( .D(n2200), .CK(clk), .RN(n1491), .Q(
        \gbuff[18][19] ) );
  DFFRX1 \gbuff_reg[18][18]  ( .D(n2201), .CK(clk), .RN(n1491), .Q(
        \gbuff[18][18] ) );
  DFFRX1 \gbuff_reg[18][17]  ( .D(n2202), .CK(clk), .RN(n1491), .Q(
        \gbuff[18][17] ) );
  DFFRX1 \gbuff_reg[18][16]  ( .D(n2203), .CK(clk), .RN(n1491), .Q(
        \gbuff[18][16] ) );
  DFFRX1 \gbuff_reg[18][15]  ( .D(n2204), .CK(clk), .RN(n1491), .Q(
        \gbuff[18][15] ) );
  DFFRX1 \gbuff_reg[18][14]  ( .D(n2205), .CK(clk), .RN(n1491), .Q(
        \gbuff[18][14] ) );
  DFFRX1 \gbuff_reg[18][13]  ( .D(n2206), .CK(clk), .RN(n1491), .Q(
        \gbuff[18][13] ) );
  DFFRX1 \gbuff_reg[18][12]  ( .D(n2207), .CK(clk), .RN(n1491), .Q(
        \gbuff[18][12] ) );
  DFFRX1 \gbuff_reg[18][11]  ( .D(n2208), .CK(clk), .RN(n1490), .Q(
        \gbuff[18][11] ) );
  DFFRX1 \gbuff_reg[18][10]  ( .D(n2209), .CK(clk), .RN(n1490), .Q(
        \gbuff[18][10] ) );
  DFFRX1 \gbuff_reg[18][9]  ( .D(n2210), .CK(clk), .RN(n1490), .Q(
        \gbuff[18][9] ) );
  DFFRX1 \gbuff_reg[18][8]  ( .D(n2211), .CK(clk), .RN(n1490), .Q(
        \gbuff[18][8] ) );
  DFFRX1 \gbuff_reg[18][7]  ( .D(n2212), .CK(clk), .RN(n1490), .Q(
        \gbuff[18][7] ) );
  DFFRX1 \gbuff_reg[18][6]  ( .D(n2213), .CK(clk), .RN(n1490), .Q(
        \gbuff[18][6] ) );
  DFFRX1 \gbuff_reg[18][5]  ( .D(n2214), .CK(clk), .RN(n1490), .Q(
        \gbuff[18][5] ) );
  DFFRX1 \gbuff_reg[18][4]  ( .D(n2215), .CK(clk), .RN(n1490), .Q(
        \gbuff[18][4] ) );
  DFFRX1 \gbuff_reg[18][3]  ( .D(n2216), .CK(clk), .RN(n1490), .Q(
        \gbuff[18][3] ) );
  DFFRX1 \gbuff_reg[18][2]  ( .D(n2217), .CK(clk), .RN(n1490), .Q(
        \gbuff[18][2] ) );
  DFFRX1 \gbuff_reg[18][1]  ( .D(n2218), .CK(clk), .RN(n1490), .Q(
        \gbuff[18][1] ) );
  DFFRX1 \gbuff_reg[18][0]  ( .D(n2219), .CK(clk), .RN(n1490), .Q(
        \gbuff[18][0] ) );
  DFFRX1 \gbuff_reg[14][31]  ( .D(n2316), .CK(clk), .RN(n1481), .Q(
        \gbuff[14][31] ) );
  DFFRX1 \gbuff_reg[14][30]  ( .D(n2317), .CK(clk), .RN(n1481), .Q(
        \gbuff[14][30] ) );
  DFFRX1 \gbuff_reg[14][29]  ( .D(n2318), .CK(clk), .RN(n1481), .Q(
        \gbuff[14][29] ) );
  DFFRX1 \gbuff_reg[14][28]  ( .D(n2319), .CK(clk), .RN(n1481), .Q(
        \gbuff[14][28] ) );
  DFFRX1 \gbuff_reg[14][27]  ( .D(n2320), .CK(clk), .RN(n1481), .Q(
        \gbuff[14][27] ) );
  DFFRX1 \gbuff_reg[14][26]  ( .D(n2321), .CK(clk), .RN(n1481), .Q(
        \gbuff[14][26] ) );
  DFFRX1 \gbuff_reg[14][25]  ( .D(n2322), .CK(clk), .RN(n1481), .Q(
        \gbuff[14][25] ) );
  DFFRX1 \gbuff_reg[14][24]  ( .D(n2323), .CK(clk), .RN(n1481), .Q(
        \gbuff[14][24] ) );
  DFFRX1 \gbuff_reg[14][23]  ( .D(n2324), .CK(clk), .RN(n1481), .Q(
        \gbuff[14][23] ) );
  DFFRX1 \gbuff_reg[14][22]  ( .D(n2325), .CK(clk), .RN(n1481), .Q(
        \gbuff[14][22] ) );
  DFFRX1 \gbuff_reg[14][21]  ( .D(n2326), .CK(clk), .RN(n1481), .Q(
        \gbuff[14][21] ) );
  DFFRX1 \gbuff_reg[14][20]  ( .D(n2327), .CK(clk), .RN(n1481), .Q(
        \gbuff[14][20] ) );
  DFFRX1 \gbuff_reg[14][19]  ( .D(n2328), .CK(clk), .RN(n1480), .Q(
        \gbuff[14][19] ) );
  DFFRX1 \gbuff_reg[14][18]  ( .D(n2329), .CK(clk), .RN(n1480), .Q(
        \gbuff[14][18] ) );
  DFFRX1 \gbuff_reg[14][17]  ( .D(n2330), .CK(clk), .RN(n1480), .Q(
        \gbuff[14][17] ) );
  DFFRX1 \gbuff_reg[14][16]  ( .D(n2331), .CK(clk), .RN(n1480), .Q(
        \gbuff[14][16] ) );
  DFFRX1 \gbuff_reg[14][15]  ( .D(n2332), .CK(clk), .RN(n1480), .Q(
        \gbuff[14][15] ) );
  DFFRX1 \gbuff_reg[14][14]  ( .D(n2333), .CK(clk), .RN(n1480), .Q(
        \gbuff[14][14] ) );
  DFFRX1 \gbuff_reg[14][13]  ( .D(n2334), .CK(clk), .RN(n1480), .Q(
        \gbuff[14][13] ) );
  DFFRX1 \gbuff_reg[14][12]  ( .D(n2335), .CK(clk), .RN(n1480), .Q(
        \gbuff[14][12] ) );
  DFFRX1 \gbuff_reg[14][11]  ( .D(n2336), .CK(clk), .RN(n1480), .Q(
        \gbuff[14][11] ) );
  DFFRX1 \gbuff_reg[14][10]  ( .D(n2337), .CK(clk), .RN(n1480), .Q(
        \gbuff[14][10] ) );
  DFFRX1 \gbuff_reg[14][9]  ( .D(n2338), .CK(clk), .RN(n1480), .Q(
        \gbuff[14][9] ) );
  DFFRX1 \gbuff_reg[14][8]  ( .D(n2339), .CK(clk), .RN(n1480), .Q(
        \gbuff[14][8] ) );
  DFFRX1 \gbuff_reg[14][7]  ( .D(n2340), .CK(clk), .RN(n1479), .Q(
        \gbuff[14][7] ) );
  DFFRX1 \gbuff_reg[14][6]  ( .D(n2341), .CK(clk), .RN(n1479), .Q(
        \gbuff[14][6] ) );
  DFFRX1 \gbuff_reg[14][5]  ( .D(n2342), .CK(clk), .RN(n1479), .Q(
        \gbuff[14][5] ) );
  DFFRX1 \gbuff_reg[14][4]  ( .D(n2343), .CK(clk), .RN(n1479), .Q(
        \gbuff[14][4] ) );
  DFFRX1 \gbuff_reg[14][3]  ( .D(n2344), .CK(clk), .RN(n1479), .Q(
        \gbuff[14][3] ) );
  DFFRX1 \gbuff_reg[14][2]  ( .D(n2345), .CK(clk), .RN(n1479), .Q(
        \gbuff[14][2] ) );
  DFFRX1 \gbuff_reg[14][1]  ( .D(n2346), .CK(clk), .RN(n1479), .Q(
        \gbuff[14][1] ) );
  DFFRX1 \gbuff_reg[14][0]  ( .D(n2347), .CK(clk), .RN(n1479), .Q(
        \gbuff[14][0] ) );
  DFFRX1 \gbuff_reg[10][31]  ( .D(n2444), .CK(clk), .RN(n1471), .Q(
        \gbuff[10][31] ) );
  DFFRX1 \gbuff_reg[10][30]  ( .D(n2445), .CK(clk), .RN(n1471), .Q(
        \gbuff[10][30] ) );
  DFFRX1 \gbuff_reg[10][29]  ( .D(n2446), .CK(clk), .RN(n1471), .Q(
        \gbuff[10][29] ) );
  DFFRX1 \gbuff_reg[10][28]  ( .D(n2447), .CK(clk), .RN(n1471), .Q(
        \gbuff[10][28] ) );
  DFFRX1 \gbuff_reg[10][27]  ( .D(n2448), .CK(clk), .RN(n1470), .Q(
        \gbuff[10][27] ) );
  DFFRX1 \gbuff_reg[10][26]  ( .D(n2449), .CK(clk), .RN(n1470), .Q(
        \gbuff[10][26] ) );
  DFFRX1 \gbuff_reg[10][25]  ( .D(n2450), .CK(clk), .RN(n1470), .Q(
        \gbuff[10][25] ) );
  DFFRX1 \gbuff_reg[10][24]  ( .D(n2451), .CK(clk), .RN(n1470), .Q(
        \gbuff[10][24] ) );
  DFFRX1 \gbuff_reg[10][23]  ( .D(n2452), .CK(clk), .RN(n1470), .Q(
        \gbuff[10][23] ) );
  DFFRX1 \gbuff_reg[10][22]  ( .D(n2453), .CK(clk), .RN(n1470), .Q(
        \gbuff[10][22] ) );
  DFFRX1 \gbuff_reg[10][21]  ( .D(n2454), .CK(clk), .RN(n1470), .Q(
        \gbuff[10][21] ) );
  DFFRX1 \gbuff_reg[10][20]  ( .D(n2455), .CK(clk), .RN(n1470), .Q(
        \gbuff[10][20] ) );
  DFFRX1 \gbuff_reg[10][19]  ( .D(n2456), .CK(clk), .RN(n1470), .Q(
        \gbuff[10][19] ) );
  DFFRX1 \gbuff_reg[10][18]  ( .D(n2457), .CK(clk), .RN(n1470), .Q(
        \gbuff[10][18] ) );
  DFFRX1 \gbuff_reg[10][17]  ( .D(n2458), .CK(clk), .RN(n1470), .Q(
        \gbuff[10][17] ) );
  DFFRX1 \gbuff_reg[10][16]  ( .D(n2459), .CK(clk), .RN(n1470), .Q(
        \gbuff[10][16] ) );
  DFFRX1 \gbuff_reg[10][15]  ( .D(n2460), .CK(clk), .RN(n1469), .Q(
        \gbuff[10][15] ) );
  DFFRX1 \gbuff_reg[10][14]  ( .D(n2461), .CK(clk), .RN(n1469), .Q(
        \gbuff[10][14] ) );
  DFFRX1 \gbuff_reg[10][13]  ( .D(n2462), .CK(clk), .RN(n1469), .Q(
        \gbuff[10][13] ) );
  DFFRX1 \gbuff_reg[10][12]  ( .D(n2463), .CK(clk), .RN(n1469), .Q(
        \gbuff[10][12] ) );
  DFFRX1 \gbuff_reg[10][11]  ( .D(n2464), .CK(clk), .RN(n1469), .Q(
        \gbuff[10][11] ) );
  DFFRX1 \gbuff_reg[10][10]  ( .D(n2465), .CK(clk), .RN(n1469), .Q(
        \gbuff[10][10] ) );
  DFFRX1 \gbuff_reg[10][9]  ( .D(n2466), .CK(clk), .RN(n1469), .Q(
        \gbuff[10][9] ) );
  DFFRX1 \gbuff_reg[10][8]  ( .D(n2467), .CK(clk), .RN(n1469), .Q(
        \gbuff[10][8] ) );
  DFFRX1 \gbuff_reg[10][7]  ( .D(n2468), .CK(clk), .RN(n1469), .Q(
        \gbuff[10][7] ) );
  DFFRX1 \gbuff_reg[10][6]  ( .D(n2469), .CK(clk), .RN(n1469), .Q(
        \gbuff[10][6] ) );
  DFFRX1 \gbuff_reg[10][5]  ( .D(n2470), .CK(clk), .RN(n1469), .Q(
        \gbuff[10][5] ) );
  DFFRX1 \gbuff_reg[10][4]  ( .D(n2471), .CK(clk), .RN(n1469), .Q(
        \gbuff[10][4] ) );
  DFFRX1 \gbuff_reg[10][3]  ( .D(n2472), .CK(clk), .RN(n1468), .Q(
        \gbuff[10][3] ) );
  DFFRX1 \gbuff_reg[10][2]  ( .D(n2473), .CK(clk), .RN(n1468), .Q(
        \gbuff[10][2] ) );
  DFFRX1 \gbuff_reg[10][1]  ( .D(n2474), .CK(clk), .RN(n1468), .Q(
        \gbuff[10][1] ) );
  DFFRX1 \gbuff_reg[10][0]  ( .D(n2475), .CK(clk), .RN(n1468), .Q(
        \gbuff[10][0] ) );
  DFFRX1 \gbuff_reg[6][31]  ( .D(n2572), .CK(clk), .RN(n1460), .Q(
        \gbuff[6][31] ) );
  DFFRX1 \gbuff_reg[6][30]  ( .D(n2573), .CK(clk), .RN(n1460), .Q(
        \gbuff[6][30] ) );
  DFFRX1 \gbuff_reg[6][29]  ( .D(n2574), .CK(clk), .RN(n1460), .Q(
        \gbuff[6][29] ) );
  DFFRX1 \gbuff_reg[6][28]  ( .D(n2575), .CK(clk), .RN(n1460), .Q(
        \gbuff[6][28] ) );
  DFFRX1 \gbuff_reg[6][27]  ( .D(n2576), .CK(clk), .RN(n1460), .Q(
        \gbuff[6][27] ) );
  DFFRX1 \gbuff_reg[6][26]  ( .D(n2577), .CK(clk), .RN(n1460), .Q(
        \gbuff[6][26] ) );
  DFFRX1 \gbuff_reg[6][25]  ( .D(n2578), .CK(clk), .RN(n1460), .Q(
        \gbuff[6][25] ) );
  DFFRX1 \gbuff_reg[6][24]  ( .D(n2579), .CK(clk), .RN(n1460), .Q(
        \gbuff[6][24] ) );
  DFFRX1 \gbuff_reg[6][23]  ( .D(n2580), .CK(clk), .RN(n1459), .Q(
        \gbuff[6][23] ) );
  DFFRX1 \gbuff_reg[6][22]  ( .D(n2581), .CK(clk), .RN(n1459), .Q(
        \gbuff[6][22] ) );
  DFFRX1 \gbuff_reg[6][21]  ( .D(n2582), .CK(clk), .RN(n1459), .Q(
        \gbuff[6][21] ) );
  DFFRX1 \gbuff_reg[6][20]  ( .D(n2583), .CK(clk), .RN(n1459), .Q(
        \gbuff[6][20] ) );
  DFFRX1 \gbuff_reg[6][19]  ( .D(n2584), .CK(clk), .RN(n1459), .Q(
        \gbuff[6][19] ) );
  DFFRX1 \gbuff_reg[6][18]  ( .D(n2585), .CK(clk), .RN(n1459), .Q(
        \gbuff[6][18] ) );
  DFFRX1 \gbuff_reg[6][17]  ( .D(n2586), .CK(clk), .RN(n1459), .Q(
        \gbuff[6][17] ) );
  DFFRX1 \gbuff_reg[6][16]  ( .D(n2587), .CK(clk), .RN(n1459), .Q(
        \gbuff[6][16] ) );
  DFFRX1 \gbuff_reg[6][15]  ( .D(n2588), .CK(clk), .RN(n1459), .Q(
        \gbuff[6][15] ) );
  DFFRX1 \gbuff_reg[6][14]  ( .D(n2589), .CK(clk), .RN(n1459), .Q(
        \gbuff[6][14] ) );
  DFFRX1 \gbuff_reg[6][13]  ( .D(n2590), .CK(clk), .RN(n1459), .Q(
        \gbuff[6][13] ) );
  DFFRX1 \gbuff_reg[6][12]  ( .D(n2591), .CK(clk), .RN(n1459), .Q(
        \gbuff[6][12] ) );
  DFFRX1 \gbuff_reg[6][11]  ( .D(n2592), .CK(clk), .RN(n1458), .Q(
        \gbuff[6][11] ) );
  DFFRX1 \gbuff_reg[6][10]  ( .D(n2593), .CK(clk), .RN(n1458), .Q(
        \gbuff[6][10] ) );
  DFFRX1 \gbuff_reg[6][9]  ( .D(n2594), .CK(clk), .RN(n1458), .Q(\gbuff[6][9] ) );
  DFFRX1 \gbuff_reg[6][8]  ( .D(n2595), .CK(clk), .RN(n1458), .Q(\gbuff[6][8] ) );
  DFFRX1 \gbuff_reg[6][7]  ( .D(n2596), .CK(clk), .RN(n1458), .Q(\gbuff[6][7] ) );
  DFFRX1 \gbuff_reg[6][6]  ( .D(n2597), .CK(clk), .RN(n1458), .Q(\gbuff[6][6] ) );
  DFFRX1 \gbuff_reg[6][5]  ( .D(n2598), .CK(clk), .RN(n1458), .Q(\gbuff[6][5] ) );
  DFFRX1 \gbuff_reg[6][4]  ( .D(n2599), .CK(clk), .RN(n1458), .Q(\gbuff[6][4] ) );
  DFFRX1 \gbuff_reg[6][3]  ( .D(n2600), .CK(clk), .RN(n1458), .Q(\gbuff[6][3] ) );
  DFFRX1 \gbuff_reg[6][2]  ( .D(n2601), .CK(clk), .RN(n1458), .Q(\gbuff[6][2] ) );
  DFFRX1 \gbuff_reg[6][1]  ( .D(n2602), .CK(clk), .RN(n1458), .Q(\gbuff[6][1] ) );
  DFFRX1 \gbuff_reg[6][0]  ( .D(n2603), .CK(clk), .RN(n1458), .Q(\gbuff[6][0] ) );
  DFFRX1 \gbuff_reg[2][31]  ( .D(n2700), .CK(clk), .RN(n1449), .Q(
        \gbuff[2][31] ) );
  DFFRX1 \gbuff_reg[2][30]  ( .D(n2701), .CK(clk), .RN(n1449), .Q(
        \gbuff[2][30] ) );
  DFFRX1 \gbuff_reg[2][29]  ( .D(n2702), .CK(clk), .RN(n1449), .Q(
        \gbuff[2][29] ) );
  DFFRX1 \gbuff_reg[2][28]  ( .D(n2703), .CK(clk), .RN(n1449), .Q(
        \gbuff[2][28] ) );
  DFFRX1 \gbuff_reg[2][27]  ( .D(n2704), .CK(clk), .RN(n1449), .Q(
        \gbuff[2][27] ) );
  DFFRX1 \gbuff_reg[2][26]  ( .D(n2705), .CK(clk), .RN(n1449), .Q(
        \gbuff[2][26] ) );
  DFFRX1 \gbuff_reg[2][25]  ( .D(n2706), .CK(clk), .RN(n1449), .Q(
        \gbuff[2][25] ) );
  DFFRX1 \gbuff_reg[2][24]  ( .D(n2707), .CK(clk), .RN(n1449), .Q(
        \gbuff[2][24] ) );
  DFFRX1 \gbuff_reg[2][23]  ( .D(n2708), .CK(clk), .RN(n1449), .Q(
        \gbuff[2][23] ) );
  DFFRX1 \gbuff_reg[2][22]  ( .D(n2709), .CK(clk), .RN(n1449), .Q(
        \gbuff[2][22] ) );
  DFFRX1 \gbuff_reg[2][21]  ( .D(n2710), .CK(clk), .RN(n1449), .Q(
        \gbuff[2][21] ) );
  DFFRX1 \gbuff_reg[2][20]  ( .D(n2711), .CK(clk), .RN(n1449), .Q(
        \gbuff[2][20] ) );
  DFFRX1 \gbuff_reg[2][19]  ( .D(n2712), .CK(clk), .RN(n1448), .Q(
        \gbuff[2][19] ) );
  DFFRX1 \gbuff_reg[2][18]  ( .D(n2713), .CK(clk), .RN(n1448), .Q(
        \gbuff[2][18] ) );
  DFFRX1 \gbuff_reg[2][17]  ( .D(n2714), .CK(clk), .RN(n1448), .Q(
        \gbuff[2][17] ) );
  DFFRX1 \gbuff_reg[2][16]  ( .D(n2715), .CK(clk), .RN(n1448), .Q(
        \gbuff[2][16] ) );
  DFFRX1 \gbuff_reg[2][15]  ( .D(n2716), .CK(clk), .RN(n1448), .Q(
        \gbuff[2][15] ) );
  DFFRX1 \gbuff_reg[2][14]  ( .D(n2717), .CK(clk), .RN(n1448), .Q(
        \gbuff[2][14] ) );
  DFFRX1 \gbuff_reg[2][13]  ( .D(n2718), .CK(clk), .RN(n1448), .Q(
        \gbuff[2][13] ) );
  DFFRX1 \gbuff_reg[2][12]  ( .D(n2719), .CK(clk), .RN(n1448), .Q(
        \gbuff[2][12] ) );
  DFFRX1 \gbuff_reg[2][11]  ( .D(n2720), .CK(clk), .RN(n1448), .Q(
        \gbuff[2][11] ) );
  DFFRX1 \gbuff_reg[2][10]  ( .D(n2721), .CK(clk), .RN(n1448), .Q(
        \gbuff[2][10] ) );
  DFFRX1 \gbuff_reg[2][9]  ( .D(n2722), .CK(clk), .RN(n1448), .Q(\gbuff[2][9] ) );
  DFFRX1 \gbuff_reg[2][8]  ( .D(n2723), .CK(clk), .RN(n1448), .Q(\gbuff[2][8] ) );
  DFFRX1 \gbuff_reg[2][7]  ( .D(n2724), .CK(clk), .RN(n1447), .Q(\gbuff[2][7] ) );
  DFFRX1 \gbuff_reg[2][6]  ( .D(n2725), .CK(clk), .RN(n1447), .Q(\gbuff[2][6] ) );
  DFFRX1 \gbuff_reg[2][5]  ( .D(n2726), .CK(clk), .RN(n1447), .Q(\gbuff[2][5] ) );
  DFFRX1 \gbuff_reg[2][4]  ( .D(n2727), .CK(clk), .RN(n1447), .Q(\gbuff[2][4] ) );
  DFFRX1 \gbuff_reg[2][3]  ( .D(n2728), .CK(clk), .RN(n1447), .Q(\gbuff[2][3] ) );
  DFFRX1 \gbuff_reg[2][2]  ( .D(n2729), .CK(clk), .RN(n1447), .Q(\gbuff[2][2] ) );
  DFFRX1 \gbuff_reg[2][1]  ( .D(n2730), .CK(clk), .RN(n1447), .Q(\gbuff[2][1] ) );
  DFFRX1 \gbuff_reg[2][0]  ( .D(n2731), .CK(clk), .RN(n1447), .Q(\gbuff[2][0] ) );
  EDFFX1 \data_out_reg[31]  ( .D(N16), .E(n1730), .CK(clk), .Q(data_out[31])
         );
  EDFFX1 \data_out_reg[30]  ( .D(N17), .E(n1729), .CK(clk), .Q(data_out[30])
         );
  EDFFX1 \data_out_reg[29]  ( .D(N18), .E(n1730), .CK(clk), .Q(data_out[29])
         );
  EDFFX1 \data_out_reg[28]  ( .D(N19), .E(n1729), .CK(clk), .Q(data_out[28])
         );
  EDFFX1 \data_out_reg[27]  ( .D(N20), .E(n1730), .CK(clk), .Q(data_out[27])
         );
  EDFFX1 \data_out_reg[26]  ( .D(N21), .E(n1729), .CK(clk), .Q(data_out[26])
         );
  EDFFX1 \data_out_reg[25]  ( .D(N22), .E(n1730), .CK(clk), .Q(data_out[25])
         );
  EDFFX1 \data_out_reg[24]  ( .D(N23), .E(n1729), .CK(clk), .Q(data_out[24])
         );
  EDFFX1 \data_out_reg[23]  ( .D(N24), .E(n1730), .CK(clk), .Q(data_out[23])
         );
  EDFFX1 \data_out_reg[22]  ( .D(N25), .E(n1730), .CK(clk), .Q(data_out[22])
         );
  EDFFX1 \data_out_reg[21]  ( .D(N26), .E(n1730), .CK(clk), .Q(data_out[21])
         );
  EDFFX1 \data_out_reg[20]  ( .D(N27), .E(n1730), .CK(clk), .Q(data_out[20])
         );
  EDFFX1 \data_out_reg[19]  ( .D(N28), .E(n1730), .CK(clk), .Q(data_out[19])
         );
  EDFFX1 \data_out_reg[18]  ( .D(N29), .E(n1730), .CK(clk), .Q(data_out[18])
         );
  EDFFX1 \data_out_reg[17]  ( .D(N30), .E(n1730), .CK(clk), .Q(data_out[17])
         );
  EDFFX1 \data_out_reg[16]  ( .D(N31), .E(n1730), .CK(clk), .Q(data_out[16])
         );
  EDFFX1 \data_out_reg[15]  ( .D(N32), .E(n1730), .CK(clk), .Q(data_out[15])
         );
  EDFFX1 \data_out_reg[14]  ( .D(N33), .E(n1730), .CK(clk), .Q(data_out[14])
         );
  EDFFX1 \data_out_reg[13]  ( .D(N34), .E(n1730), .CK(clk), .Q(data_out[13])
         );
  EDFFX1 \data_out_reg[12]  ( .D(N35), .E(n1730), .CK(clk), .Q(data_out[12])
         );
  EDFFX1 \data_out_reg[11]  ( .D(N36), .E(n1729), .CK(clk), .Q(data_out[11])
         );
  EDFFX1 \data_out_reg[10]  ( .D(N37), .E(n1729), .CK(clk), .Q(data_out[10])
         );
  EDFFX1 \data_out_reg[9]  ( .D(N38), .E(n1729), .CK(clk), .Q(data_out[9]) );
  EDFFX1 \data_out_reg[8]  ( .D(N39), .E(n1729), .CK(clk), .Q(data_out[8]) );
  EDFFX1 \data_out_reg[7]  ( .D(N40), .E(n1729), .CK(clk), .Q(data_out[7]) );
  EDFFX1 \data_out_reg[6]  ( .D(N41), .E(n1729), .CK(clk), .Q(data_out[6]) );
  EDFFX1 \data_out_reg[5]  ( .D(N42), .E(n1729), .CK(clk), .Q(data_out[5]) );
  EDFFX1 \data_out_reg[4]  ( .D(N43), .E(n1729), .CK(clk), .Q(data_out[4]) );
  EDFFX1 \data_out_reg[3]  ( .D(N44), .E(n1729), .CK(clk), .Q(data_out[3]) );
  EDFFX1 \data_out_reg[2]  ( .D(N45), .E(n1729), .CK(clk), .Q(data_out[2]) );
  EDFFX1 \data_out_reg[1]  ( .D(N46), .E(n1729), .CK(clk), .Q(data_out[1]) );
  EDFFX1 \data_out_reg[0]  ( .D(N47), .E(n1729), .CK(clk), .Q(data_out[0]) );
  NOR4BX1 U2 ( .AN(wr_en), .B(index[5]), .C(index[7]), .D(index[6]), .Y(n2815)
         );
  NOR3BX2 U3 ( .AN(n2815), .B(n1736), .C(n1738), .Y(n2823) );
  NOR3BX2 U4 ( .AN(n2815), .B(n1738), .C(n1737), .Y(n2814) );
  NAND2X1 U5 ( .A(n2824), .B(n2823), .Y(n1) );
  NAND2X1 U6 ( .A(n2820), .B(n2823), .Y(n2) );
  NAND2X1 U7 ( .A(n2818), .B(n2823), .Y(n3) );
  NAND2X1 U8 ( .A(n2817), .B(n2823), .Y(n4) );
  NAND2X1 U9 ( .A(n2816), .B(n2823), .Y(n5) );
  NAND2X1 U10 ( .A(n2814), .B(n2820), .Y(n6) );
  NAND2X1 U11 ( .A(n2814), .B(n2818), .Y(n7) );
  NAND2X1 U12 ( .A(n2814), .B(n2817), .Y(n8) );
  NAND2X1 U13 ( .A(n2814), .B(n2816), .Y(n9) );
  NAND2X1 U14 ( .A(n2814), .B(n2824), .Y(n10) );
  NAND2X1 U15 ( .A(n2814), .B(n2822), .Y(n11) );
  NAND2X1 U16 ( .A(n2814), .B(n2819), .Y(n12) );
  NAND2X1 U17 ( .A(n2814), .B(n2821), .Y(n13) );
  NAND2X1 U18 ( .A(n2822), .B(n2823), .Y(n14) );
  NAND2X1 U19 ( .A(n2821), .B(n2823), .Y(n15) );
  NAND2X1 U20 ( .A(n2819), .B(n2823), .Y(n16) );
  CLKINVX1 U21 ( .A(n1732), .Y(n1731) );
  CLKINVX1 U22 ( .A(n1734), .Y(n1733) );
  NOR3X1 U23 ( .A(n1733), .B(n1735), .C(n1731), .Y(n2824) );
  NOR3X1 U24 ( .A(n1733), .B(n1735), .C(n1732), .Y(n2822) );
  NOR3X1 U25 ( .A(n1731), .B(n1735), .C(n1734), .Y(n2821) );
  NOR3X1 U26 ( .A(n1732), .B(n1735), .C(n1734), .Y(n2820) );
  NOR2X1 U27 ( .A(wr_en), .B(rst), .Y(N81) );
  CLKINVX1 U28 ( .A(N11), .Y(n1734) );
  CLKINVX1 U29 ( .A(N10), .Y(n1732) );
  CLKINVX1 U30 ( .A(N13), .Y(n1737) );
  CLKINVX1 U31 ( .A(data_in[0]), .Y(n1771) );
  CLKINVX1 U32 ( .A(data_in[1]), .Y(n1770) );
  CLKINVX1 U33 ( .A(data_in[2]), .Y(n1769) );
  CLKINVX1 U34 ( .A(data_in[3]), .Y(n1768) );
  CLKINVX1 U35 ( .A(data_in[4]), .Y(n1767) );
  CLKINVX1 U36 ( .A(data_in[5]), .Y(n1766) );
  CLKINVX1 U37 ( .A(data_in[6]), .Y(n1765) );
  CLKINVX1 U38 ( .A(data_in[7]), .Y(n1764) );
  CLKINVX1 U39 ( .A(data_in[8]), .Y(n1763) );
  CLKINVX1 U40 ( .A(data_in[9]), .Y(n1762) );
  CLKINVX1 U41 ( .A(data_in[10]), .Y(n1761) );
  CLKINVX1 U42 ( .A(data_in[11]), .Y(n1760) );
  CLKINVX1 U43 ( .A(data_in[12]), .Y(n1759) );
  CLKINVX1 U44 ( .A(data_in[13]), .Y(n1758) );
  CLKINVX1 U45 ( .A(data_in[14]), .Y(n1757) );
  CLKINVX1 U46 ( .A(data_in[15]), .Y(n1756) );
  CLKINVX1 U47 ( .A(data_in[16]), .Y(n1755) );
  CLKINVX1 U48 ( .A(data_in[17]), .Y(n1754) );
  CLKINVX1 U49 ( .A(data_in[18]), .Y(n1753) );
  CLKINVX1 U50 ( .A(data_in[19]), .Y(n1752) );
  CLKINVX1 U51 ( .A(data_in[20]), .Y(n1751) );
  CLKINVX1 U52 ( .A(data_in[21]), .Y(n1750) );
  CLKINVX1 U53 ( .A(data_in[22]), .Y(n1749) );
  CLKINVX1 U54 ( .A(data_in[23]), .Y(n1748) );
  CLKINVX1 U55 ( .A(data_in[24]), .Y(n1747) );
  CLKINVX1 U56 ( .A(data_in[25]), .Y(n1746) );
  CLKINVX1 U57 ( .A(data_in[26]), .Y(n1745) );
  CLKINVX1 U58 ( .A(data_in[27]), .Y(n1744) );
  CLKINVX1 U59 ( .A(data_in[28]), .Y(n1743) );
  CLKINVX1 U60 ( .A(data_in[29]), .Y(n1742) );
  CLKINVX1 U61 ( .A(data_in[30]), .Y(n1741) );
  CLKINVX1 U62 ( .A(data_in[31]), .Y(n1740) );
  CLKINVX1 U63 ( .A(rst), .Y(n1739) );
  CLKBUFX3 U64 ( .A(n1436), .Y(n1419) );
  CLKBUFX3 U65 ( .A(n1436), .Y(n1420) );
  CLKBUFX3 U66 ( .A(n1436), .Y(n1421) );
  CLKBUFX3 U67 ( .A(n1437), .Y(n1422) );
  CLKBUFX3 U68 ( .A(n1437), .Y(n1423) );
  CLKBUFX3 U69 ( .A(n1437), .Y(n1424) );
  CLKBUFX3 U70 ( .A(n1437), .Y(n1425) );
  CLKBUFX3 U71 ( .A(n1417), .Y(n1426) );
  CLKBUFX3 U72 ( .A(n1417), .Y(n1427) );
  CLKBUFX3 U73 ( .A(n1437), .Y(n1428) );
  CLKBUFX3 U74 ( .A(n1437), .Y(n1429) );
  CLKBUFX3 U75 ( .A(n1417), .Y(n1430) );
  CLKBUFX3 U76 ( .A(n1417), .Y(n1431) );
  CLKBUFX3 U77 ( .A(n1436), .Y(n1432) );
  CLKBUFX3 U78 ( .A(n1417), .Y(n1433) );
  CLKBUFX3 U79 ( .A(n1417), .Y(n1434) );
  CLKBUFX3 U80 ( .A(n1417), .Y(n1435) );
  CLKBUFX3 U81 ( .A(n1404), .Y(n1400) );
  CLKBUFX3 U82 ( .A(N11), .Y(n1401) );
  CLKBUFX3 U83 ( .A(n1398), .Y(n1402) );
  CLKBUFX3 U84 ( .A(n1401), .Y(n1403) );
  CLKBUFX3 U85 ( .A(n1401), .Y(n1404) );
  CLKBUFX3 U86 ( .A(n1398), .Y(n1405) );
  CLKBUFX3 U87 ( .A(n1401), .Y(n1406) );
  CLKBUFX3 U88 ( .A(n1416), .Y(n1407) );
  CLKBUFX3 U89 ( .A(n1398), .Y(n1408) );
  CLKBUFX3 U90 ( .A(n1398), .Y(n1409) );
  CLKBUFX3 U91 ( .A(n1406), .Y(n1410) );
  CLKBUFX3 U92 ( .A(n1401), .Y(n1411) );
  CLKBUFX3 U93 ( .A(n1398), .Y(n1412) );
  CLKBUFX3 U94 ( .A(n1403), .Y(n1413) );
  CLKBUFX3 U95 ( .A(n1398), .Y(n1414) );
  CLKBUFX3 U96 ( .A(n1398), .Y(n1415) );
  CLKBUFX3 U97 ( .A(n1401), .Y(n1416) );
  CLKBUFX3 U98 ( .A(n1436), .Y(n1418) );
  CLKBUFX3 U99 ( .A(n1), .Y(n1728) );
  CLKBUFX3 U100 ( .A(n1), .Y(n1727) );
  CLKBUFX3 U101 ( .A(n10), .Y(n1703) );
  CLKBUFX3 U102 ( .A(n11), .Y(n1700) );
  CLKBUFX3 U103 ( .A(n12), .Y(n1691) );
  CLKBUFX3 U104 ( .A(n2799), .Y(n1643) );
  CLKBUFX3 U105 ( .A(n2798), .Y(n1640) );
  CLKBUFX3 U106 ( .A(n2797), .Y(n1637) );
  CLKBUFX3 U107 ( .A(n2796), .Y(n1634) );
  CLKBUFX3 U108 ( .A(n1), .Y(n1726) );
  CLKBUFX3 U109 ( .A(n14), .Y(n1725) );
  CLKBUFX3 U110 ( .A(n15), .Y(n1722) );
  CLKBUFX3 U111 ( .A(n16), .Y(n1716) );
  CLKBUFX3 U112 ( .A(n10), .Y(n1704) );
  CLKBUFX3 U113 ( .A(n11), .Y(n1701) );
  CLKBUFX3 U114 ( .A(n13), .Y(n1698) );
  CLKBUFX3 U115 ( .A(n6), .Y(n1695) );
  CLKBUFX3 U116 ( .A(n12), .Y(n1692) );
  CLKBUFX3 U117 ( .A(n7), .Y(n1689) );
  CLKBUFX3 U118 ( .A(n8), .Y(n1686) );
  CLKBUFX3 U119 ( .A(n9), .Y(n1683) );
  CLKBUFX3 U120 ( .A(n14), .Y(n1723) );
  CLKBUFX3 U121 ( .A(n14), .Y(n1724) );
  CLKBUFX3 U122 ( .A(n15), .Y(n1720) );
  CLKBUFX3 U123 ( .A(n15), .Y(n1721) );
  CLKBUFX3 U124 ( .A(n1717), .Y(n1718) );
  CLKBUFX3 U125 ( .A(n1717), .Y(n1719) );
  CLKBUFX3 U126 ( .A(n16), .Y(n1714) );
  CLKBUFX3 U127 ( .A(n16), .Y(n1715) );
  CLKBUFX3 U128 ( .A(n1711), .Y(n1712) );
  CLKBUFX3 U129 ( .A(n1711), .Y(n1713) );
  CLKBUFX3 U130 ( .A(n1708), .Y(n1709) );
  CLKBUFX3 U131 ( .A(n1708), .Y(n1710) );
  CLKBUFX3 U132 ( .A(n1705), .Y(n1706) );
  CLKBUFX3 U133 ( .A(n1705), .Y(n1707) );
  CLKBUFX3 U134 ( .A(n10), .Y(n1702) );
  CLKBUFX3 U135 ( .A(n11), .Y(n1699) );
  CLKBUFX3 U136 ( .A(n13), .Y(n1696) );
  CLKBUFX3 U137 ( .A(n13), .Y(n1697) );
  CLKBUFX3 U138 ( .A(n1693), .Y(n1694) );
  CLKBUFX3 U139 ( .A(n12), .Y(n1690) );
  CLKBUFX3 U140 ( .A(n1687), .Y(n1688) );
  CLKBUFX3 U141 ( .A(n1684), .Y(n1685) );
  CLKBUFX3 U142 ( .A(n1681), .Y(n1682) );
  CLKBUFX3 U143 ( .A(n1678), .Y(n1679) );
  CLKBUFX3 U144 ( .A(n1675), .Y(n1676) );
  CLKBUFX3 U145 ( .A(n1672), .Y(n1673) );
  CLKBUFX3 U146 ( .A(n1669), .Y(n1670) );
  CLKBUFX3 U147 ( .A(n1666), .Y(n1667) );
  CLKBUFX3 U148 ( .A(n2807), .Y(n1663) );
  CLKBUFX3 U149 ( .A(n2807), .Y(n1664) );
  CLKBUFX3 U150 ( .A(n2806), .Y(n1660) );
  CLKBUFX3 U151 ( .A(n2806), .Y(n1661) );
  CLKBUFX3 U152 ( .A(n2805), .Y(n1657) );
  CLKBUFX3 U153 ( .A(n2805), .Y(n1658) );
  CLKBUFX3 U154 ( .A(n1654), .Y(n1655) );
  CLKBUFX3 U155 ( .A(n1651), .Y(n1652) );
  CLKBUFX3 U156 ( .A(n1648), .Y(n1649) );
  CLKBUFX3 U157 ( .A(n1645), .Y(n1646) );
  CLKBUFX3 U158 ( .A(n2799), .Y(n1642) );
  CLKBUFX3 U159 ( .A(n2798), .Y(n1639) );
  CLKBUFX3 U160 ( .A(n2797), .Y(n1636) );
  CLKBUFX3 U161 ( .A(n2796), .Y(n1633) );
  CLKBUFX3 U162 ( .A(n1398), .Y(n1399) );
  CLKBUFX3 U163 ( .A(N11), .Y(n1398) );
  CLKBUFX3 U164 ( .A(n1678), .Y(n1680) );
  CLKBUFX3 U165 ( .A(n1675), .Y(n1677) );
  CLKBUFX3 U166 ( .A(n1672), .Y(n1674) );
  CLKBUFX3 U167 ( .A(n1669), .Y(n1671) );
  CLKBUFX3 U168 ( .A(n1666), .Y(n1668) );
  CLKBUFX3 U169 ( .A(n2807), .Y(n1665) );
  CLKBUFX3 U170 ( .A(n2806), .Y(n1662) );
  CLKBUFX3 U171 ( .A(n2805), .Y(n1659) );
  CLKBUFX3 U172 ( .A(n1654), .Y(n1656) );
  CLKBUFX3 U173 ( .A(n1651), .Y(n1653) );
  CLKBUFX3 U174 ( .A(n1648), .Y(n1650) );
  CLKBUFX3 U175 ( .A(n1645), .Y(n1647) );
  CLKBUFX3 U176 ( .A(n2799), .Y(n1644) );
  CLKBUFX3 U177 ( .A(n2798), .Y(n1641) );
  CLKBUFX3 U178 ( .A(n2797), .Y(n1638) );
  CLKBUFX3 U179 ( .A(n2796), .Y(n1635) );
  CLKBUFX3 U180 ( .A(n1736), .Y(n1391) );
  CLKBUFX3 U181 ( .A(N13), .Y(n1392) );
  CLKBUFX3 U182 ( .A(N13), .Y(n1393) );
  CLKBUFX3 U183 ( .A(N13), .Y(n1394) );
  CLKBUFX3 U184 ( .A(n1557), .Y(n1442) );
  CLKBUFX3 U185 ( .A(n1557), .Y(n1443) );
  CLKBUFX3 U186 ( .A(n1556), .Y(n1444) );
  CLKBUFX3 U187 ( .A(n1556), .Y(n1445) );
  CLKBUFX3 U188 ( .A(n1555), .Y(n1446) );
  CLKBUFX3 U189 ( .A(n1555), .Y(n1447) );
  CLKBUFX3 U190 ( .A(n1554), .Y(n1448) );
  CLKBUFX3 U191 ( .A(n1554), .Y(n1449) );
  CLKBUFX3 U192 ( .A(n1553), .Y(n1450) );
  CLKBUFX3 U193 ( .A(n1553), .Y(n1451) );
  CLKBUFX3 U194 ( .A(n1552), .Y(n1452) );
  CLKBUFX3 U195 ( .A(n1552), .Y(n1453) );
  CLKBUFX3 U196 ( .A(n1551), .Y(n1454) );
  CLKBUFX3 U197 ( .A(n1551), .Y(n1455) );
  CLKBUFX3 U198 ( .A(n1550), .Y(n1456) );
  CLKBUFX3 U199 ( .A(n1550), .Y(n1457) );
  CLKBUFX3 U200 ( .A(n1549), .Y(n1458) );
  CLKBUFX3 U201 ( .A(n1549), .Y(n1459) );
  CLKBUFX3 U202 ( .A(n1548), .Y(n1460) );
  CLKBUFX3 U203 ( .A(n1548), .Y(n1461) );
  CLKBUFX3 U204 ( .A(n1547), .Y(n1462) );
  CLKBUFX3 U205 ( .A(n1547), .Y(n1463) );
  CLKBUFX3 U206 ( .A(n1546), .Y(n1464) );
  CLKBUFX3 U207 ( .A(n1546), .Y(n1465) );
  CLKBUFX3 U208 ( .A(n1545), .Y(n1466) );
  CLKBUFX3 U209 ( .A(n1545), .Y(n1467) );
  CLKBUFX3 U210 ( .A(n1544), .Y(n1468) );
  CLKBUFX3 U211 ( .A(n1544), .Y(n1469) );
  CLKBUFX3 U212 ( .A(n1543), .Y(n1470) );
  CLKBUFX3 U213 ( .A(n1543), .Y(n1471) );
  CLKBUFX3 U214 ( .A(n1542), .Y(n1472) );
  CLKBUFX3 U215 ( .A(n1542), .Y(n1473) );
  CLKBUFX3 U216 ( .A(n1541), .Y(n1474) );
  CLKBUFX3 U217 ( .A(n1541), .Y(n1475) );
  CLKBUFX3 U218 ( .A(n1540), .Y(n1476) );
  CLKBUFX3 U219 ( .A(n1540), .Y(n1477) );
  CLKBUFX3 U220 ( .A(n1539), .Y(n1478) );
  CLKBUFX3 U221 ( .A(n1539), .Y(n1479) );
  CLKBUFX3 U222 ( .A(n1538), .Y(n1480) );
  CLKBUFX3 U223 ( .A(n1538), .Y(n1481) );
  CLKBUFX3 U224 ( .A(n1537), .Y(n1482) );
  CLKBUFX3 U225 ( .A(n1537), .Y(n1483) );
  CLKBUFX3 U226 ( .A(n1536), .Y(n1484) );
  CLKBUFX3 U227 ( .A(n1536), .Y(n1485) );
  CLKBUFX3 U228 ( .A(n1535), .Y(n1486) );
  CLKBUFX3 U229 ( .A(n1535), .Y(n1487) );
  CLKBUFX3 U230 ( .A(n1534), .Y(n1488) );
  CLKBUFX3 U231 ( .A(n1534), .Y(n1489) );
  CLKBUFX3 U232 ( .A(n1533), .Y(n1490) );
  CLKBUFX3 U233 ( .A(n1533), .Y(n1491) );
  CLKBUFX3 U234 ( .A(n1532), .Y(n1492) );
  CLKBUFX3 U235 ( .A(n1532), .Y(n1493) );
  CLKBUFX3 U236 ( .A(n1531), .Y(n1494) );
  CLKBUFX3 U237 ( .A(n1531), .Y(n1495) );
  CLKBUFX3 U238 ( .A(n1530), .Y(n1496) );
  CLKBUFX3 U239 ( .A(n1530), .Y(n1497) );
  CLKBUFX3 U240 ( .A(n1565), .Y(n1498) );
  CLKBUFX3 U241 ( .A(n1543), .Y(n1499) );
  CLKBUFX3 U242 ( .A(n1545), .Y(n1500) );
  CLKBUFX3 U243 ( .A(n1544), .Y(n1501) );
  CLKBUFX3 U244 ( .A(n1529), .Y(n1502) );
  CLKBUFX3 U245 ( .A(n1529), .Y(n1503) );
  CLKBUFX3 U246 ( .A(n1528), .Y(n1504) );
  CLKBUFX3 U247 ( .A(n1528), .Y(n1505) );
  CLKBUFX3 U248 ( .A(n1566), .Y(n1506) );
  CLKBUFX3 U249 ( .A(n1547), .Y(n1507) );
  CLKBUFX3 U250 ( .A(n1566), .Y(n1508) );
  CLKBUFX3 U251 ( .A(n1548), .Y(n1509) );
  CLKBUFX3 U252 ( .A(n1550), .Y(n1510) );
  CLKBUFX3 U253 ( .A(n1549), .Y(n1511) );
  CLKBUFX3 U254 ( .A(n1566), .Y(n1512) );
  CLKBUFX3 U255 ( .A(n1546), .Y(n1513) );
  CLKBUFX3 U256 ( .A(n1567), .Y(n1514) );
  CLKBUFX3 U257 ( .A(n1551), .Y(n1515) );
  CLKBUFX3 U258 ( .A(n1567), .Y(n1516) );
  CLKBUFX3 U259 ( .A(n1552), .Y(n1517) );
  CLKBUFX3 U260 ( .A(n1567), .Y(n1518) );
  CLKBUFX3 U261 ( .A(n1553), .Y(n1519) );
  CLKBUFX3 U262 ( .A(n1555), .Y(n1520) );
  CLKBUFX3 U263 ( .A(n1554), .Y(n1521) );
  CLKBUFX3 U264 ( .A(n1568), .Y(n1522) );
  CLKBUFX3 U265 ( .A(n1556), .Y(n1523) );
  CLKBUFX3 U266 ( .A(n1568), .Y(n1524) );
  CLKBUFX3 U267 ( .A(n1557), .Y(n1525) );
  CLKBUFX3 U268 ( .A(n1568), .Y(n1526) );
  CLKBUFX3 U269 ( .A(n1441), .Y(n1527) );
  CLKBUFX3 U270 ( .A(n2813), .Y(n1678) );
  CLKBUFX3 U271 ( .A(n2811), .Y(n1675) );
  CLKBUFX3 U272 ( .A(n2810), .Y(n1672) );
  CLKBUFX3 U273 ( .A(n2809), .Y(n1669) );
  CLKBUFX3 U274 ( .A(n2808), .Y(n1666) );
  CLKBUFX3 U275 ( .A(n2804), .Y(n1654) );
  CLKBUFX3 U276 ( .A(n2802), .Y(n1651) );
  CLKBUFX3 U277 ( .A(n2801), .Y(n1648) );
  CLKBUFX3 U278 ( .A(n2800), .Y(n1645) );
  CLKBUFX3 U279 ( .A(n2), .Y(n1717) );
  CLKBUFX3 U280 ( .A(n3), .Y(n1711) );
  CLKBUFX3 U281 ( .A(n4), .Y(n1708) );
  CLKBUFX3 U282 ( .A(n5), .Y(n1705) );
  CLKBUFX3 U283 ( .A(n6), .Y(n1693) );
  CLKBUFX3 U284 ( .A(n7), .Y(n1687) );
  CLKBUFX3 U285 ( .A(n8), .Y(n1684) );
  CLKBUFX3 U286 ( .A(n9), .Y(n1681) );
  CLKBUFX3 U287 ( .A(n1437), .Y(n1417) );
  CLKBUFX3 U288 ( .A(n1735), .Y(n1395) );
  CLKBUFX3 U289 ( .A(N12), .Y(n1396) );
  CLKBUFX3 U290 ( .A(n1735), .Y(n1397) );
  CLKBUFX3 U291 ( .A(n1558), .Y(n1557) );
  CLKBUFX3 U292 ( .A(n1558), .Y(n1556) );
  CLKBUFX3 U293 ( .A(n1558), .Y(n1555) );
  CLKBUFX3 U294 ( .A(n1558), .Y(n1554) );
  CLKBUFX3 U295 ( .A(n1559), .Y(n1553) );
  CLKBUFX3 U296 ( .A(n1559), .Y(n1552) );
  CLKBUFX3 U297 ( .A(n1559), .Y(n1551) );
  CLKBUFX3 U298 ( .A(n1559), .Y(n1550) );
  CLKBUFX3 U299 ( .A(n1560), .Y(n1549) );
  CLKBUFX3 U300 ( .A(n1560), .Y(n1548) );
  CLKBUFX3 U301 ( .A(n1560), .Y(n1547) );
  CLKBUFX3 U302 ( .A(n1560), .Y(n1546) );
  CLKBUFX3 U303 ( .A(n1561), .Y(n1545) );
  CLKBUFX3 U304 ( .A(n1561), .Y(n1544) );
  CLKBUFX3 U305 ( .A(n1561), .Y(n1543) );
  CLKBUFX3 U306 ( .A(n1561), .Y(n1542) );
  CLKBUFX3 U307 ( .A(n1562), .Y(n1541) );
  CLKBUFX3 U308 ( .A(n1562), .Y(n1540) );
  CLKBUFX3 U309 ( .A(n1562), .Y(n1539) );
  CLKBUFX3 U310 ( .A(n1562), .Y(n1538) );
  CLKBUFX3 U311 ( .A(n1563), .Y(n1537) );
  CLKBUFX3 U312 ( .A(n1563), .Y(n1536) );
  CLKBUFX3 U313 ( .A(n1563), .Y(n1535) );
  CLKBUFX3 U314 ( .A(n1563), .Y(n1534) );
  CLKBUFX3 U315 ( .A(n1564), .Y(n1533) );
  CLKBUFX3 U316 ( .A(n1564), .Y(n1532) );
  CLKBUFX3 U317 ( .A(n1564), .Y(n1531) );
  CLKBUFX3 U318 ( .A(n1564), .Y(n1530) );
  CLKBUFX3 U319 ( .A(n1565), .Y(n1529) );
  CLKBUFX3 U320 ( .A(n1565), .Y(n1528) );
  NAND2X1 U321 ( .A(n2812), .B(n2824), .Y(n2813) );
  NAND2X1 U322 ( .A(n2812), .B(n2822), .Y(n2811) );
  NAND2X1 U323 ( .A(n2812), .B(n2821), .Y(n2810) );
  NAND2X1 U324 ( .A(n2812), .B(n2820), .Y(n2809) );
  NAND2X1 U325 ( .A(n2803), .B(n2824), .Y(n2804) );
  NAND2X1 U326 ( .A(n2803), .B(n2822), .Y(n2802) );
  NAND2X1 U327 ( .A(n2803), .B(n2821), .Y(n2801) );
  NAND2X1 U328 ( .A(n2803), .B(n2820), .Y(n2800) );
  NAND2X1 U329 ( .A(n2812), .B(n2819), .Y(n2808) );
  NAND2X1 U330 ( .A(n2812), .B(n2818), .Y(n2807) );
  NAND2X1 U331 ( .A(n2812), .B(n2817), .Y(n2806) );
  NAND2X1 U332 ( .A(n2812), .B(n2816), .Y(n2805) );
  NAND2X1 U333 ( .A(n2803), .B(n2819), .Y(n2799) );
  NAND2X1 U334 ( .A(n2803), .B(n2818), .Y(n2798) );
  NAND2X1 U335 ( .A(n2803), .B(n2817), .Y(n2797) );
  NAND2X1 U336 ( .A(n2803), .B(n2816), .Y(n2796) );
  CLKBUFX3 U337 ( .A(n1731), .Y(n1436) );
  CLKBUFX3 U338 ( .A(n1731), .Y(n1437) );
  CLKBUFX3 U339 ( .A(n1738), .Y(n1390) );
  CLKBUFX3 U340 ( .A(n1438), .Y(n1558) );
  CLKBUFX3 U341 ( .A(n1438), .Y(n1559) );
  CLKBUFX3 U342 ( .A(n1438), .Y(n1560) );
  CLKBUFX3 U343 ( .A(n1439), .Y(n1561) );
  CLKBUFX3 U344 ( .A(n1439), .Y(n1562) );
  CLKBUFX3 U345 ( .A(n1439), .Y(n1563) );
  CLKBUFX3 U346 ( .A(n1440), .Y(n1564) );
  CLKBUFX3 U347 ( .A(n1440), .Y(n1565) );
  CLKBUFX3 U348 ( .A(n1440), .Y(n1566) );
  CLKBUFX3 U349 ( .A(n1441), .Y(n1567) );
  CLKBUFX3 U350 ( .A(n1441), .Y(n1568) );
  CLKBUFX3 U351 ( .A(N81), .Y(n1729) );
  CLKBUFX3 U352 ( .A(N81), .Y(n1730) );
  AND3X2 U353 ( .A(n2815), .B(n1737), .C(n1738), .Y(n2812) );
  AND3X2 U354 ( .A(n1736), .B(n2815), .C(n1738), .Y(n2803) );
  AND3X2 U355 ( .A(n1735), .B(n1732), .C(n1734), .Y(n2819) );
  AND3X2 U356 ( .A(n1735), .B(n1731), .C(n1734), .Y(n2818) );
  AND3X2 U357 ( .A(n1735), .B(n1733), .C(n1732), .Y(n2817) );
  AND3X2 U358 ( .A(n1735), .B(n1733), .C(n1731), .Y(n2816) );
  CLKBUFX3 U359 ( .A(n1771), .Y(n1632) );
  CLKBUFX3 U360 ( .A(n1770), .Y(n1630) );
  CLKBUFX3 U361 ( .A(n1769), .Y(n1628) );
  CLKBUFX3 U362 ( .A(n1768), .Y(n1626) );
  CLKBUFX3 U363 ( .A(n1767), .Y(n1624) );
  CLKBUFX3 U364 ( .A(n1766), .Y(n1622) );
  CLKBUFX3 U365 ( .A(n1765), .Y(n1620) );
  CLKBUFX3 U366 ( .A(n1764), .Y(n1618) );
  CLKBUFX3 U367 ( .A(n1763), .Y(n1616) );
  CLKBUFX3 U368 ( .A(n1762), .Y(n1614) );
  CLKBUFX3 U369 ( .A(n1761), .Y(n1612) );
  CLKBUFX3 U370 ( .A(n1760), .Y(n1610) );
  CLKBUFX3 U371 ( .A(n1759), .Y(n1608) );
  CLKBUFX3 U372 ( .A(n1758), .Y(n1606) );
  CLKBUFX3 U373 ( .A(n1757), .Y(n1604) );
  CLKBUFX3 U374 ( .A(n1756), .Y(n1602) );
  CLKBUFX3 U375 ( .A(n1755), .Y(n1600) );
  CLKBUFX3 U376 ( .A(n1754), .Y(n1598) );
  CLKBUFX3 U377 ( .A(n1753), .Y(n1596) );
  CLKBUFX3 U378 ( .A(n1752), .Y(n1594) );
  CLKBUFX3 U379 ( .A(n1751), .Y(n1592) );
  CLKBUFX3 U380 ( .A(n1750), .Y(n1590) );
  CLKBUFX3 U381 ( .A(n1749), .Y(n1588) );
  CLKBUFX3 U382 ( .A(n1748), .Y(n1586) );
  CLKBUFX3 U383 ( .A(n1771), .Y(n1631) );
  CLKBUFX3 U384 ( .A(n1770), .Y(n1629) );
  CLKBUFX3 U385 ( .A(n1769), .Y(n1627) );
  CLKBUFX3 U386 ( .A(n1768), .Y(n1625) );
  CLKBUFX3 U387 ( .A(n1767), .Y(n1623) );
  CLKBUFX3 U388 ( .A(n1766), .Y(n1621) );
  CLKBUFX3 U389 ( .A(n1765), .Y(n1619) );
  CLKBUFX3 U390 ( .A(n1764), .Y(n1617) );
  CLKBUFX3 U391 ( .A(n1763), .Y(n1615) );
  CLKBUFX3 U392 ( .A(n1762), .Y(n1613) );
  CLKBUFX3 U393 ( .A(n1761), .Y(n1611) );
  CLKBUFX3 U394 ( .A(n1760), .Y(n1609) );
  CLKBUFX3 U395 ( .A(n1759), .Y(n1607) );
  CLKBUFX3 U396 ( .A(n1758), .Y(n1605) );
  CLKBUFX3 U397 ( .A(n1757), .Y(n1603) );
  CLKBUFX3 U398 ( .A(n1756), .Y(n1601) );
  CLKBUFX3 U399 ( .A(n1755), .Y(n1599) );
  CLKBUFX3 U400 ( .A(n1754), .Y(n1597) );
  CLKBUFX3 U401 ( .A(n1753), .Y(n1595) );
  CLKBUFX3 U402 ( .A(n1752), .Y(n1593) );
  CLKBUFX3 U403 ( .A(n1751), .Y(n1591) );
  CLKBUFX3 U404 ( .A(n1750), .Y(n1589) );
  CLKBUFX3 U405 ( .A(n1749), .Y(n1587) );
  CLKBUFX3 U406 ( .A(n1748), .Y(n1585) );
  CLKINVX1 U407 ( .A(n1737), .Y(n1736) );
  CLKBUFX3 U408 ( .A(n1747), .Y(n1584) );
  CLKBUFX3 U409 ( .A(n1746), .Y(n1582) );
  CLKBUFX3 U410 ( .A(n1745), .Y(n1580) );
  CLKBUFX3 U411 ( .A(n1744), .Y(n1578) );
  CLKBUFX3 U412 ( .A(n1743), .Y(n1576) );
  CLKBUFX3 U413 ( .A(n1742), .Y(n1574) );
  CLKBUFX3 U414 ( .A(n1741), .Y(n1572) );
  CLKBUFX3 U415 ( .A(n1740), .Y(n1570) );
  CLKBUFX3 U416 ( .A(n1747), .Y(n1583) );
  CLKBUFX3 U417 ( .A(n1746), .Y(n1581) );
  CLKBUFX3 U418 ( .A(n1745), .Y(n1579) );
  CLKBUFX3 U419 ( .A(n1744), .Y(n1577) );
  CLKBUFX3 U420 ( .A(n1743), .Y(n1575) );
  CLKBUFX3 U421 ( .A(n1742), .Y(n1573) );
  CLKBUFX3 U422 ( .A(n1741), .Y(n1571) );
  CLKBUFX3 U423 ( .A(n1740), .Y(n1569) );
  CLKBUFX3 U424 ( .A(n1739), .Y(n1438) );
  CLKBUFX3 U425 ( .A(n1739), .Y(n1439) );
  CLKBUFX3 U426 ( .A(n1739), .Y(n1440) );
  CLKBUFX3 U427 ( .A(n1739), .Y(n1441) );
  OAI2BB2XL U428 ( .B0(n1727), .B1(n1748), .A0N(\gbuff[0][23] ), .A1N(n1727), 
        .Y(n2772) );
  OAI2BB2XL U429 ( .B0(n1727), .B1(n1746), .A0N(\gbuff[0][25] ), .A1N(n1728), 
        .Y(n2770) );
  OAI2BB2XL U430 ( .B0(n1727), .B1(n1745), .A0N(\gbuff[0][26] ), .A1N(n1728), 
        .Y(n2769) );
  OAI2BB2XL U431 ( .B0(n1727), .B1(n1744), .A0N(\gbuff[0][27] ), .A1N(n1728), 
        .Y(n2768) );
  OAI2BB2XL U432 ( .B0(n1727), .B1(n1743), .A0N(\gbuff[0][28] ), .A1N(n1728), 
        .Y(n2767) );
  OAI2BB2XL U433 ( .B0(n1727), .B1(n1742), .A0N(\gbuff[0][29] ), .A1N(n1728), 
        .Y(n2766) );
  OAI2BB2XL U434 ( .B0(n1727), .B1(n1741), .A0N(\gbuff[0][30] ), .A1N(n1726), 
        .Y(n2765) );
  OAI2BB2XL U435 ( .B0(n1727), .B1(n1740), .A0N(\gbuff[0][31] ), .A1N(n1728), 
        .Y(n2764) );
  OAI2BB2XL U436 ( .B0(n1586), .B1(n1723), .A0N(\gbuff[1][23] ), .A1N(n1724), 
        .Y(n2740) );
  OAI2BB2XL U437 ( .B0(n1582), .B1(n1724), .A0N(\gbuff[1][25] ), .A1N(n1725), 
        .Y(n2738) );
  OAI2BB2XL U438 ( .B0(n1580), .B1(n1723), .A0N(\gbuff[1][26] ), .A1N(n1725), 
        .Y(n2737) );
  OAI2BB2XL U439 ( .B0(n1578), .B1(n1724), .A0N(\gbuff[1][27] ), .A1N(n1725), 
        .Y(n2736) );
  OAI2BB2XL U440 ( .B0(n1576), .B1(n1723), .A0N(\gbuff[1][28] ), .A1N(n1725), 
        .Y(n2735) );
  OAI2BB2XL U441 ( .B0(n1574), .B1(n1724), .A0N(\gbuff[1][29] ), .A1N(n1725), 
        .Y(n2734) );
  OAI2BB2XL U442 ( .B0(n1572), .B1(n14), .A0N(\gbuff[1][30] ), .A1N(n1723), 
        .Y(n2733) );
  OAI2BB2XL U443 ( .B0(n1570), .B1(n14), .A0N(\gbuff[1][31] ), .A1N(n1724), 
        .Y(n2732) );
  OAI2BB2XL U444 ( .B0(n1585), .B1(n1720), .A0N(\gbuff[2][23] ), .A1N(n1721), 
        .Y(n2708) );
  OAI2BB2XL U445 ( .B0(n1581), .B1(n1721), .A0N(\gbuff[2][25] ), .A1N(n1722), 
        .Y(n2706) );
  OAI2BB2XL U446 ( .B0(n1579), .B1(n1720), .A0N(\gbuff[2][26] ), .A1N(n1722), 
        .Y(n2705) );
  OAI2BB2XL U447 ( .B0(n1577), .B1(n1721), .A0N(\gbuff[2][27] ), .A1N(n1722), 
        .Y(n2704) );
  OAI2BB2XL U448 ( .B0(n1575), .B1(n1720), .A0N(\gbuff[2][28] ), .A1N(n1722), 
        .Y(n2703) );
  OAI2BB2XL U449 ( .B0(n1573), .B1(n1721), .A0N(\gbuff[2][29] ), .A1N(n1722), 
        .Y(n2702) );
  OAI2BB2XL U450 ( .B0(n1571), .B1(n15), .A0N(\gbuff[2][30] ), .A1N(n1720), 
        .Y(n2701) );
  OAI2BB2XL U451 ( .B0(n1569), .B1(n15), .A0N(\gbuff[2][31] ), .A1N(n1721), 
        .Y(n2700) );
  OAI2BB2XL U452 ( .B0(n1586), .B1(n1717), .A0N(\gbuff[3][23] ), .A1N(n2), .Y(
        n2676) );
  OAI2BB2XL U453 ( .B0(n1582), .B1(n1717), .A0N(\gbuff[3][25] ), .A1N(n1717), 
        .Y(n2674) );
  OAI2BB2XL U454 ( .B0(n1580), .B1(n2), .A0N(\gbuff[3][26] ), .A1N(n1717), .Y(
        n2673) );
  OAI2BB2XL U455 ( .B0(n1578), .B1(n1717), .A0N(\gbuff[3][27] ), .A1N(n1718), 
        .Y(n2672) );
  OAI2BB2XL U456 ( .B0(n1576), .B1(n1717), .A0N(\gbuff[3][28] ), .A1N(n1719), 
        .Y(n2671) );
  OAI2BB2XL U457 ( .B0(n1574), .B1(n2), .A0N(\gbuff[3][29] ), .A1N(n1717), .Y(
        n2670) );
  OAI2BB2XL U458 ( .B0(n1572), .B1(n2), .A0N(\gbuff[3][30] ), .A1N(n1718), .Y(
        n2669) );
  OAI2BB2XL U459 ( .B0(n1570), .B1(n2), .A0N(\gbuff[3][31] ), .A1N(n1719), .Y(
        n2668) );
  OAI2BB2XL U460 ( .B0(n1585), .B1(n1714), .A0N(\gbuff[4][23] ), .A1N(n16), 
        .Y(n2644) );
  OAI2BB2XL U461 ( .B0(n1581), .B1(n1715), .A0N(\gbuff[4][25] ), .A1N(n1716), 
        .Y(n2642) );
  OAI2BB2XL U462 ( .B0(n1579), .B1(n1714), .A0N(\gbuff[4][26] ), .A1N(n1716), 
        .Y(n2641) );
  OAI2BB2XL U463 ( .B0(n1577), .B1(n1715), .A0N(\gbuff[4][27] ), .A1N(n1716), 
        .Y(n2640) );
  OAI2BB2XL U464 ( .B0(n1575), .B1(n1714), .A0N(\gbuff[4][28] ), .A1N(n1716), 
        .Y(n2639) );
  OAI2BB2XL U465 ( .B0(n1573), .B1(n1715), .A0N(\gbuff[4][29] ), .A1N(n1716), 
        .Y(n2638) );
  OAI2BB2XL U466 ( .B0(n1571), .B1(n1714), .A0N(\gbuff[4][30] ), .A1N(n1714), 
        .Y(n2637) );
  OAI2BB2XL U467 ( .B0(n1569), .B1(n1715), .A0N(\gbuff[4][31] ), .A1N(n1715), 
        .Y(n2636) );
  OAI2BB2XL U468 ( .B0(n1748), .B1(n1711), .A0N(\gbuff[5][23] ), .A1N(n3), .Y(
        n2612) );
  OAI2BB2XL U469 ( .B0(n1746), .B1(n1711), .A0N(\gbuff[5][25] ), .A1N(n1711), 
        .Y(n2610) );
  OAI2BB2XL U470 ( .B0(n1745), .B1(n3), .A0N(\gbuff[5][26] ), .A1N(n1711), .Y(
        n2609) );
  OAI2BB2XL U471 ( .B0(n1744), .B1(n1711), .A0N(\gbuff[5][27] ), .A1N(n1712), 
        .Y(n2608) );
  OAI2BB2XL U472 ( .B0(n1743), .B1(n1711), .A0N(\gbuff[5][28] ), .A1N(n1713), 
        .Y(n2607) );
  OAI2BB2XL U473 ( .B0(n1742), .B1(n3), .A0N(\gbuff[5][29] ), .A1N(n1711), .Y(
        n2606) );
  OAI2BB2XL U474 ( .B0(n1741), .B1(n3), .A0N(\gbuff[5][30] ), .A1N(n1712), .Y(
        n2605) );
  OAI2BB2XL U475 ( .B0(n1740), .B1(n3), .A0N(\gbuff[5][31] ), .A1N(n1713), .Y(
        n2604) );
  OAI2BB2XL U476 ( .B0(n1748), .B1(n1708), .A0N(\gbuff[6][23] ), .A1N(n4), .Y(
        n2580) );
  OAI2BB2XL U477 ( .B0(n1746), .B1(n1708), .A0N(\gbuff[6][25] ), .A1N(n1708), 
        .Y(n2578) );
  OAI2BB2XL U478 ( .B0(n1745), .B1(n4), .A0N(\gbuff[6][26] ), .A1N(n1708), .Y(
        n2577) );
  OAI2BB2XL U479 ( .B0(n1744), .B1(n1708), .A0N(\gbuff[6][27] ), .A1N(n1709), 
        .Y(n2576) );
  OAI2BB2XL U480 ( .B0(n1743), .B1(n1708), .A0N(\gbuff[6][28] ), .A1N(n1710), 
        .Y(n2575) );
  OAI2BB2XL U481 ( .B0(n1742), .B1(n4), .A0N(\gbuff[6][29] ), .A1N(n1708), .Y(
        n2574) );
  OAI2BB2XL U482 ( .B0(n1741), .B1(n4), .A0N(\gbuff[6][30] ), .A1N(n1709), .Y(
        n2573) );
  OAI2BB2XL U483 ( .B0(n1740), .B1(n4), .A0N(\gbuff[6][31] ), .A1N(n1710), .Y(
        n2572) );
  OAI2BB2XL U484 ( .B0(n1748), .B1(n1705), .A0N(\gbuff[7][23] ), .A1N(n5), .Y(
        n2548) );
  OAI2BB2XL U485 ( .B0(n1746), .B1(n1705), .A0N(\gbuff[7][25] ), .A1N(n1705), 
        .Y(n2546) );
  OAI2BB2XL U486 ( .B0(n1745), .B1(n5), .A0N(\gbuff[7][26] ), .A1N(n1705), .Y(
        n2545) );
  OAI2BB2XL U487 ( .B0(n1744), .B1(n1705), .A0N(\gbuff[7][27] ), .A1N(n1706), 
        .Y(n2544) );
  OAI2BB2XL U488 ( .B0(n1743), .B1(n1705), .A0N(\gbuff[7][28] ), .A1N(n1707), 
        .Y(n2543) );
  OAI2BB2XL U489 ( .B0(n1742), .B1(n5), .A0N(\gbuff[7][29] ), .A1N(n1705), .Y(
        n2542) );
  OAI2BB2XL U490 ( .B0(n1741), .B1(n5), .A0N(\gbuff[7][30] ), .A1N(n1706), .Y(
        n2541) );
  OAI2BB2XL U491 ( .B0(n1740), .B1(n5), .A0N(\gbuff[7][31] ), .A1N(n1707), .Y(
        n2540) );
  OAI2BB2XL U492 ( .B0(n1586), .B1(n1703), .A0N(\gbuff[8][23] ), .A1N(n1703), 
        .Y(n2516) );
  OAI2BB2XL U493 ( .B0(n1582), .B1(n1703), .A0N(\gbuff[8][25] ), .A1N(n1704), 
        .Y(n2514) );
  OAI2BB2XL U494 ( .B0(n1580), .B1(n1703), .A0N(\gbuff[8][26] ), .A1N(n1704), 
        .Y(n2513) );
  OAI2BB2XL U495 ( .B0(n1578), .B1(n1703), .A0N(\gbuff[8][27] ), .A1N(n1704), 
        .Y(n2512) );
  OAI2BB2XL U496 ( .B0(n1576), .B1(n1703), .A0N(\gbuff[8][28] ), .A1N(n1704), 
        .Y(n2511) );
  OAI2BB2XL U497 ( .B0(n1574), .B1(n1703), .A0N(\gbuff[8][29] ), .A1N(n1704), 
        .Y(n2510) );
  OAI2BB2XL U498 ( .B0(n1572), .B1(n1703), .A0N(\gbuff[8][30] ), .A1N(n1702), 
        .Y(n2509) );
  OAI2BB2XL U499 ( .B0(n1570), .B1(n1703), .A0N(\gbuff[8][31] ), .A1N(n1704), 
        .Y(n2508) );
  OAI2BB2XL U500 ( .B0(n1586), .B1(n1700), .A0N(\gbuff[9][23] ), .A1N(n1700), 
        .Y(n2484) );
  OAI2BB2XL U501 ( .B0(n1582), .B1(n1700), .A0N(\gbuff[9][25] ), .A1N(n1701), 
        .Y(n2482) );
  OAI2BB2XL U502 ( .B0(n1580), .B1(n1700), .A0N(\gbuff[9][26] ), .A1N(n1701), 
        .Y(n2481) );
  OAI2BB2XL U503 ( .B0(n1578), .B1(n1700), .A0N(\gbuff[9][27] ), .A1N(n1701), 
        .Y(n2480) );
  OAI2BB2XL U504 ( .B0(n1576), .B1(n1700), .A0N(\gbuff[9][28] ), .A1N(n1701), 
        .Y(n2479) );
  OAI2BB2XL U505 ( .B0(n1574), .B1(n1700), .A0N(\gbuff[9][29] ), .A1N(n1701), 
        .Y(n2478) );
  OAI2BB2XL U506 ( .B0(n1572), .B1(n1700), .A0N(\gbuff[9][30] ), .A1N(n1699), 
        .Y(n2477) );
  OAI2BB2XL U507 ( .B0(n1570), .B1(n1700), .A0N(\gbuff[9][31] ), .A1N(n1701), 
        .Y(n2476) );
  OAI2BB2XL U508 ( .B0(n1586), .B1(n1696), .A0N(\gbuff[10][23] ), .A1N(n1697), 
        .Y(n2452) );
  OAI2BB2XL U509 ( .B0(n1582), .B1(n1697), .A0N(\gbuff[10][25] ), .A1N(n1698), 
        .Y(n2450) );
  OAI2BB2XL U510 ( .B0(n1580), .B1(n1696), .A0N(\gbuff[10][26] ), .A1N(n1698), 
        .Y(n2449) );
  OAI2BB2XL U511 ( .B0(n1578), .B1(n1697), .A0N(\gbuff[10][27] ), .A1N(n1698), 
        .Y(n2448) );
  OAI2BB2XL U512 ( .B0(n1576), .B1(n1696), .A0N(\gbuff[10][28] ), .A1N(n1698), 
        .Y(n2447) );
  OAI2BB2XL U513 ( .B0(n1574), .B1(n1697), .A0N(\gbuff[10][29] ), .A1N(n1698), 
        .Y(n2446) );
  OAI2BB2XL U514 ( .B0(n1572), .B1(n13), .A0N(\gbuff[10][30] ), .A1N(n1696), 
        .Y(n2445) );
  OAI2BB2XL U515 ( .B0(n1570), .B1(n13), .A0N(\gbuff[10][31] ), .A1N(n1697), 
        .Y(n2444) );
  OAI2BB2XL U516 ( .B0(n1586), .B1(n1695), .A0N(\gbuff[11][23] ), .A1N(n6), 
        .Y(n2420) );
  OAI2BB2XL U517 ( .B0(n1582), .B1(n1695), .A0N(\gbuff[11][25] ), .A1N(n1695), 
        .Y(n2418) );
  OAI2BB2XL U518 ( .B0(n1580), .B1(n1695), .A0N(\gbuff[11][26] ), .A1N(n1695), 
        .Y(n2417) );
  OAI2BB2XL U519 ( .B0(n1578), .B1(n1693), .A0N(\gbuff[11][27] ), .A1N(n1695), 
        .Y(n2416) );
  OAI2BB2XL U520 ( .B0(n1576), .B1(n1693), .A0N(\gbuff[11][28] ), .A1N(n1695), 
        .Y(n2415) );
  OAI2BB2XL U521 ( .B0(n1574), .B1(n6), .A0N(\gbuff[11][29] ), .A1N(n1695), 
        .Y(n2414) );
  OAI2BB2XL U522 ( .B0(n1572), .B1(n6), .A0N(\gbuff[11][30] ), .A1N(n1694), 
        .Y(n2413) );
  OAI2BB2XL U523 ( .B0(n1570), .B1(n6), .A0N(\gbuff[11][31] ), .A1N(n1694), 
        .Y(n2412) );
  OAI2BB2XL U524 ( .B0(n1586), .B1(n1691), .A0N(\gbuff[12][23] ), .A1N(n1691), 
        .Y(n2388) );
  OAI2BB2XL U525 ( .B0(n1582), .B1(n1691), .A0N(\gbuff[12][25] ), .A1N(n1692), 
        .Y(n2386) );
  OAI2BB2XL U526 ( .B0(n1580), .B1(n1691), .A0N(\gbuff[12][26] ), .A1N(n1692), 
        .Y(n2385) );
  OAI2BB2XL U527 ( .B0(n1578), .B1(n1691), .A0N(\gbuff[12][27] ), .A1N(n1692), 
        .Y(n2384) );
  OAI2BB2XL U528 ( .B0(n1576), .B1(n1691), .A0N(\gbuff[12][28] ), .A1N(n1692), 
        .Y(n2383) );
  OAI2BB2XL U529 ( .B0(n1574), .B1(n1691), .A0N(\gbuff[12][29] ), .A1N(n1692), 
        .Y(n2382) );
  OAI2BB2XL U530 ( .B0(n1572), .B1(n1691), .A0N(\gbuff[12][30] ), .A1N(n1690), 
        .Y(n2381) );
  OAI2BB2XL U531 ( .B0(n1570), .B1(n1691), .A0N(\gbuff[12][31] ), .A1N(n1692), 
        .Y(n2380) );
  OAI2BB2XL U532 ( .B0(n1586), .B1(n1689), .A0N(\gbuff[13][23] ), .A1N(n7), 
        .Y(n2356) );
  OAI2BB2XL U533 ( .B0(n1582), .B1(n1689), .A0N(\gbuff[13][25] ), .A1N(n1689), 
        .Y(n2354) );
  OAI2BB2XL U534 ( .B0(n1580), .B1(n1689), .A0N(\gbuff[13][26] ), .A1N(n1689), 
        .Y(n2353) );
  OAI2BB2XL U535 ( .B0(n1578), .B1(n1687), .A0N(\gbuff[13][27] ), .A1N(n1689), 
        .Y(n2352) );
  OAI2BB2XL U536 ( .B0(n1576), .B1(n1687), .A0N(\gbuff[13][28] ), .A1N(n1689), 
        .Y(n2351) );
  OAI2BB2XL U537 ( .B0(n1574), .B1(n7), .A0N(\gbuff[13][29] ), .A1N(n1689), 
        .Y(n2350) );
  OAI2BB2XL U538 ( .B0(n1572), .B1(n7), .A0N(\gbuff[13][30] ), .A1N(n1688), 
        .Y(n2349) );
  OAI2BB2XL U539 ( .B0(n1570), .B1(n7), .A0N(\gbuff[13][31] ), .A1N(n1688), 
        .Y(n2348) );
  OAI2BB2XL U540 ( .B0(n1586), .B1(n1686), .A0N(\gbuff[14][23] ), .A1N(n8), 
        .Y(n2324) );
  OAI2BB2XL U541 ( .B0(n1582), .B1(n1686), .A0N(\gbuff[14][25] ), .A1N(n1686), 
        .Y(n2322) );
  OAI2BB2XL U542 ( .B0(n1580), .B1(n1686), .A0N(\gbuff[14][26] ), .A1N(n1686), 
        .Y(n2321) );
  OAI2BB2XL U543 ( .B0(n1578), .B1(n1684), .A0N(\gbuff[14][27] ), .A1N(n1686), 
        .Y(n2320) );
  OAI2BB2XL U544 ( .B0(n1576), .B1(n1684), .A0N(\gbuff[14][28] ), .A1N(n1686), 
        .Y(n2319) );
  OAI2BB2XL U545 ( .B0(n1574), .B1(n8), .A0N(\gbuff[14][29] ), .A1N(n1686), 
        .Y(n2318) );
  OAI2BB2XL U546 ( .B0(n1572), .B1(n8), .A0N(\gbuff[14][30] ), .A1N(n1685), 
        .Y(n2317) );
  OAI2BB2XL U547 ( .B0(n1570), .B1(n8), .A0N(\gbuff[14][31] ), .A1N(n1685), 
        .Y(n2316) );
  OAI2BB2XL U548 ( .B0(n1586), .B1(n1683), .A0N(\gbuff[15][23] ), .A1N(n9), 
        .Y(n2292) );
  OAI2BB2XL U549 ( .B0(n1582), .B1(n1683), .A0N(\gbuff[15][25] ), .A1N(n1683), 
        .Y(n2290) );
  OAI2BB2XL U550 ( .B0(n1580), .B1(n1683), .A0N(\gbuff[15][26] ), .A1N(n1683), 
        .Y(n2289) );
  OAI2BB2XL U551 ( .B0(n1578), .B1(n1681), .A0N(\gbuff[15][27] ), .A1N(n1683), 
        .Y(n2288) );
  OAI2BB2XL U552 ( .B0(n1576), .B1(n1681), .A0N(\gbuff[15][28] ), .A1N(n1683), 
        .Y(n2287) );
  OAI2BB2XL U553 ( .B0(n1574), .B1(n9), .A0N(\gbuff[15][29] ), .A1N(n1683), 
        .Y(n2286) );
  OAI2BB2XL U554 ( .B0(n1572), .B1(n9), .A0N(\gbuff[15][30] ), .A1N(n1682), 
        .Y(n2285) );
  OAI2BB2XL U555 ( .B0(n1570), .B1(n9), .A0N(\gbuff[15][31] ), .A1N(n1682), 
        .Y(n2284) );
  OAI2BB2XL U556 ( .B0(n1586), .B1(n1678), .A0N(\gbuff[16][23] ), .A1N(n1678), 
        .Y(n2260) );
  OAI2BB2XL U557 ( .B0(n1582), .B1(n1678), .A0N(\gbuff[16][25] ), .A1N(n1680), 
        .Y(n2258) );
  OAI2BB2XL U558 ( .B0(n1580), .B1(n2813), .A0N(\gbuff[16][26] ), .A1N(n1680), 
        .Y(n2257) );
  OAI2BB2XL U559 ( .B0(n1578), .B1(n1678), .A0N(\gbuff[16][27] ), .A1N(n1680), 
        .Y(n2256) );
  OAI2BB2XL U560 ( .B0(n1576), .B1(n1678), .A0N(\gbuff[16][28] ), .A1N(n1680), 
        .Y(n2255) );
  OAI2BB2XL U561 ( .B0(n1574), .B1(n1678), .A0N(\gbuff[16][29] ), .A1N(n1680), 
        .Y(n2254) );
  OAI2BB2XL U562 ( .B0(n1572), .B1(n1678), .A0N(\gbuff[16][30] ), .A1N(n1679), 
        .Y(n2253) );
  OAI2BB2XL U563 ( .B0(n1570), .B1(n1678), .A0N(\gbuff[16][31] ), .A1N(n2813), 
        .Y(n2252) );
  OAI2BB2XL U564 ( .B0(n1586), .B1(n1675), .A0N(\gbuff[17][23] ), .A1N(n1675), 
        .Y(n2228) );
  OAI2BB2XL U565 ( .B0(n1582), .B1(n1675), .A0N(\gbuff[17][25] ), .A1N(n1677), 
        .Y(n2226) );
  OAI2BB2XL U566 ( .B0(n1580), .B1(n2811), .A0N(\gbuff[17][26] ), .A1N(n1677), 
        .Y(n2225) );
  OAI2BB2XL U567 ( .B0(n1578), .B1(n1675), .A0N(\gbuff[17][27] ), .A1N(n1677), 
        .Y(n2224) );
  OAI2BB2XL U568 ( .B0(n1576), .B1(n1675), .A0N(\gbuff[17][28] ), .A1N(n1677), 
        .Y(n2223) );
  OAI2BB2XL U569 ( .B0(n1574), .B1(n1675), .A0N(\gbuff[17][29] ), .A1N(n1677), 
        .Y(n2222) );
  OAI2BB2XL U570 ( .B0(n1572), .B1(n1675), .A0N(\gbuff[17][30] ), .A1N(n1676), 
        .Y(n2221) );
  OAI2BB2XL U571 ( .B0(n1570), .B1(n1675), .A0N(\gbuff[17][31] ), .A1N(n2811), 
        .Y(n2220) );
  OAI2BB2XL U572 ( .B0(n1586), .B1(n1672), .A0N(\gbuff[18][23] ), .A1N(n1672), 
        .Y(n2196) );
  OAI2BB2XL U573 ( .B0(n1582), .B1(n1672), .A0N(\gbuff[18][25] ), .A1N(n1674), 
        .Y(n2194) );
  OAI2BB2XL U574 ( .B0(n1580), .B1(n2810), .A0N(\gbuff[18][26] ), .A1N(n1674), 
        .Y(n2193) );
  OAI2BB2XL U575 ( .B0(n1578), .B1(n1672), .A0N(\gbuff[18][27] ), .A1N(n1674), 
        .Y(n2192) );
  OAI2BB2XL U576 ( .B0(n1576), .B1(n1672), .A0N(\gbuff[18][28] ), .A1N(n1674), 
        .Y(n2191) );
  OAI2BB2XL U577 ( .B0(n1574), .B1(n1672), .A0N(\gbuff[18][29] ), .A1N(n1674), 
        .Y(n2190) );
  OAI2BB2XL U578 ( .B0(n1572), .B1(n1672), .A0N(\gbuff[18][30] ), .A1N(n1673), 
        .Y(n2189) );
  OAI2BB2XL U579 ( .B0(n1570), .B1(n1672), .A0N(\gbuff[18][31] ), .A1N(n2810), 
        .Y(n2188) );
  OAI2BB2XL U580 ( .B0(n1586), .B1(n1669), .A0N(\gbuff[19][23] ), .A1N(n1669), 
        .Y(n2164) );
  OAI2BB2XL U581 ( .B0(n1582), .B1(n1669), .A0N(\gbuff[19][25] ), .A1N(n1671), 
        .Y(n2162) );
  OAI2BB2XL U582 ( .B0(n1580), .B1(n2809), .A0N(\gbuff[19][26] ), .A1N(n1671), 
        .Y(n2161) );
  OAI2BB2XL U583 ( .B0(n1578), .B1(n1669), .A0N(\gbuff[19][27] ), .A1N(n1671), 
        .Y(n2160) );
  OAI2BB2XL U584 ( .B0(n1576), .B1(n1669), .A0N(\gbuff[19][28] ), .A1N(n1671), 
        .Y(n2159) );
  OAI2BB2XL U585 ( .B0(n1574), .B1(n1669), .A0N(\gbuff[19][29] ), .A1N(n1671), 
        .Y(n2158) );
  OAI2BB2XL U586 ( .B0(n1572), .B1(n1669), .A0N(\gbuff[19][30] ), .A1N(n1670), 
        .Y(n2157) );
  OAI2BB2XL U587 ( .B0(n1570), .B1(n1669), .A0N(\gbuff[19][31] ), .A1N(n2809), 
        .Y(n2156) );
  OAI2BB2XL U588 ( .B0(n1585), .B1(n2808), .A0N(\gbuff[20][23] ), .A1N(n1666), 
        .Y(n2132) );
  OAI2BB2XL U589 ( .B0(n1581), .B1(n1666), .A0N(\gbuff[20][25] ), .A1N(n1668), 
        .Y(n2130) );
  OAI2BB2XL U590 ( .B0(n1579), .B1(n1666), .A0N(\gbuff[20][26] ), .A1N(n1668), 
        .Y(n2129) );
  OAI2BB2XL U591 ( .B0(n1577), .B1(n1666), .A0N(\gbuff[20][27] ), .A1N(n1668), 
        .Y(n2128) );
  OAI2BB2XL U592 ( .B0(n1575), .B1(n1666), .A0N(\gbuff[20][28] ), .A1N(n1668), 
        .Y(n2127) );
  OAI2BB2XL U593 ( .B0(n1573), .B1(n1666), .A0N(\gbuff[20][29] ), .A1N(n1668), 
        .Y(n2126) );
  OAI2BB2XL U594 ( .B0(n1571), .B1(n1666), .A0N(\gbuff[20][30] ), .A1N(n1667), 
        .Y(n2125) );
  OAI2BB2XL U595 ( .B0(n1569), .B1(n1666), .A0N(\gbuff[20][31] ), .A1N(n1666), 
        .Y(n2124) );
  OAI2BB2XL U596 ( .B0(n1585), .B1(n1663), .A0N(\gbuff[21][23] ), .A1N(n1664), 
        .Y(n2100) );
  OAI2BB2XL U597 ( .B0(n1581), .B1(n1664), .A0N(\gbuff[21][25] ), .A1N(n1665), 
        .Y(n2098) );
  OAI2BB2XL U598 ( .B0(n1579), .B1(n1663), .A0N(\gbuff[21][26] ), .A1N(n1665), 
        .Y(n2097) );
  OAI2BB2XL U599 ( .B0(n1577), .B1(n1664), .A0N(\gbuff[21][27] ), .A1N(n1665), 
        .Y(n2096) );
  OAI2BB2XL U600 ( .B0(n1575), .B1(n2807), .A0N(\gbuff[21][28] ), .A1N(n1665), 
        .Y(n2095) );
  OAI2BB2XL U601 ( .B0(n1573), .B1(n2807), .A0N(\gbuff[21][29] ), .A1N(n1665), 
        .Y(n2094) );
  OAI2BB2XL U602 ( .B0(n1571), .B1(n2807), .A0N(\gbuff[21][30] ), .A1N(n1663), 
        .Y(n2093) );
  OAI2BB2XL U603 ( .B0(n1569), .B1(n2807), .A0N(\gbuff[21][31] ), .A1N(n1664), 
        .Y(n2092) );
  OAI2BB2XL U604 ( .B0(n1585), .B1(n1660), .A0N(\gbuff[22][23] ), .A1N(n1661), 
        .Y(n2068) );
  OAI2BB2XL U605 ( .B0(n1581), .B1(n1661), .A0N(\gbuff[22][25] ), .A1N(n1662), 
        .Y(n2066) );
  OAI2BB2XL U606 ( .B0(n1579), .B1(n1660), .A0N(\gbuff[22][26] ), .A1N(n1662), 
        .Y(n2065) );
  OAI2BB2XL U607 ( .B0(n1577), .B1(n1661), .A0N(\gbuff[22][27] ), .A1N(n1662), 
        .Y(n2064) );
  OAI2BB2XL U608 ( .B0(n1575), .B1(n2806), .A0N(\gbuff[22][28] ), .A1N(n1662), 
        .Y(n2063) );
  OAI2BB2XL U609 ( .B0(n1573), .B1(n2806), .A0N(\gbuff[22][29] ), .A1N(n1662), 
        .Y(n2062) );
  OAI2BB2XL U610 ( .B0(n1571), .B1(n2806), .A0N(\gbuff[22][30] ), .A1N(n1660), 
        .Y(n2061) );
  OAI2BB2XL U611 ( .B0(n1569), .B1(n2806), .A0N(\gbuff[22][31] ), .A1N(n1661), 
        .Y(n2060) );
  OAI2BB2XL U612 ( .B0(n1585), .B1(n1657), .A0N(\gbuff[23][23] ), .A1N(n1658), 
        .Y(n2036) );
  OAI2BB2XL U613 ( .B0(n1581), .B1(n1658), .A0N(\gbuff[23][25] ), .A1N(n1659), 
        .Y(n2034) );
  OAI2BB2XL U614 ( .B0(n1579), .B1(n1657), .A0N(\gbuff[23][26] ), .A1N(n1659), 
        .Y(n2033) );
  OAI2BB2XL U615 ( .B0(n1577), .B1(n1658), .A0N(\gbuff[23][27] ), .A1N(n1659), 
        .Y(n2032) );
  OAI2BB2XL U616 ( .B0(n1575), .B1(n2805), .A0N(\gbuff[23][28] ), .A1N(n1659), 
        .Y(n2031) );
  OAI2BB2XL U617 ( .B0(n1573), .B1(n2805), .A0N(\gbuff[23][29] ), .A1N(n1659), 
        .Y(n2030) );
  OAI2BB2XL U618 ( .B0(n1571), .B1(n2805), .A0N(\gbuff[23][30] ), .A1N(n1657), 
        .Y(n2029) );
  OAI2BB2XL U619 ( .B0(n1569), .B1(n2805), .A0N(\gbuff[23][31] ), .A1N(n1658), 
        .Y(n2028) );
  OAI2BB2XL U620 ( .B0(n1585), .B1(n1654), .A0N(\gbuff[24][23] ), .A1N(n1654), 
        .Y(n2004) );
  OAI2BB2XL U621 ( .B0(n1581), .B1(n1654), .A0N(\gbuff[24][25] ), .A1N(n1656), 
        .Y(n2002) );
  OAI2BB2XL U622 ( .B0(n1579), .B1(n2804), .A0N(\gbuff[24][26] ), .A1N(n1656), 
        .Y(n2001) );
  OAI2BB2XL U623 ( .B0(n1577), .B1(n1654), .A0N(\gbuff[24][27] ), .A1N(n1656), 
        .Y(n2000) );
  OAI2BB2XL U624 ( .B0(n1575), .B1(n1654), .A0N(\gbuff[24][28] ), .A1N(n1656), 
        .Y(n1999) );
  OAI2BB2XL U625 ( .B0(n1573), .B1(n1654), .A0N(\gbuff[24][29] ), .A1N(n1656), 
        .Y(n1998) );
  OAI2BB2XL U626 ( .B0(n1571), .B1(n1654), .A0N(\gbuff[24][30] ), .A1N(n1655), 
        .Y(n1997) );
  OAI2BB2XL U627 ( .B0(n1569), .B1(n1654), .A0N(\gbuff[24][31] ), .A1N(n2804), 
        .Y(n1996) );
  OAI2BB2XL U628 ( .B0(n1585), .B1(n1651), .A0N(\gbuff[25][23] ), .A1N(n1651), 
        .Y(n1972) );
  OAI2BB2XL U629 ( .B0(n1581), .B1(n1651), .A0N(\gbuff[25][25] ), .A1N(n1653), 
        .Y(n1970) );
  OAI2BB2XL U630 ( .B0(n1579), .B1(n2802), .A0N(\gbuff[25][26] ), .A1N(n1653), 
        .Y(n1969) );
  OAI2BB2XL U631 ( .B0(n1577), .B1(n1651), .A0N(\gbuff[25][27] ), .A1N(n1653), 
        .Y(n1968) );
  OAI2BB2XL U632 ( .B0(n1575), .B1(n1651), .A0N(\gbuff[25][28] ), .A1N(n1653), 
        .Y(n1967) );
  OAI2BB2XL U633 ( .B0(n1573), .B1(n1651), .A0N(\gbuff[25][29] ), .A1N(n1653), 
        .Y(n1966) );
  OAI2BB2XL U634 ( .B0(n1571), .B1(n1651), .A0N(\gbuff[25][30] ), .A1N(n1652), 
        .Y(n1965) );
  OAI2BB2XL U635 ( .B0(n1569), .B1(n1651), .A0N(\gbuff[25][31] ), .A1N(n2802), 
        .Y(n1964) );
  OAI2BB2XL U636 ( .B0(n1585), .B1(n1648), .A0N(\gbuff[26][23] ), .A1N(n1648), 
        .Y(n1940) );
  OAI2BB2XL U637 ( .B0(n1581), .B1(n1648), .A0N(\gbuff[26][25] ), .A1N(n1650), 
        .Y(n1938) );
  OAI2BB2XL U638 ( .B0(n1579), .B1(n2801), .A0N(\gbuff[26][26] ), .A1N(n1650), 
        .Y(n1937) );
  OAI2BB2XL U639 ( .B0(n1577), .B1(n1648), .A0N(\gbuff[26][27] ), .A1N(n1650), 
        .Y(n1936) );
  OAI2BB2XL U640 ( .B0(n1575), .B1(n1648), .A0N(\gbuff[26][28] ), .A1N(n1650), 
        .Y(n1935) );
  OAI2BB2XL U641 ( .B0(n1573), .B1(n1648), .A0N(\gbuff[26][29] ), .A1N(n1650), 
        .Y(n1934) );
  OAI2BB2XL U642 ( .B0(n1571), .B1(n1648), .A0N(\gbuff[26][30] ), .A1N(n1649), 
        .Y(n1933) );
  OAI2BB2XL U643 ( .B0(n1569), .B1(n1648), .A0N(\gbuff[26][31] ), .A1N(n2801), 
        .Y(n1932) );
  OAI2BB2XL U644 ( .B0(n1585), .B1(n1645), .A0N(\gbuff[27][23] ), .A1N(n1647), 
        .Y(n1908) );
  OAI2BB2XL U645 ( .B0(n1581), .B1(n1645), .A0N(\gbuff[27][25] ), .A1N(n1647), 
        .Y(n1906) );
  OAI2BB2XL U646 ( .B0(n1579), .B1(n1645), .A0N(\gbuff[27][26] ), .A1N(n1647), 
        .Y(n1905) );
  OAI2BB2XL U647 ( .B0(n1577), .B1(n1645), .A0N(\gbuff[27][27] ), .A1N(n1647), 
        .Y(n1904) );
  OAI2BB2XL U648 ( .B0(n1575), .B1(n1645), .A0N(\gbuff[27][28] ), .A1N(n1647), 
        .Y(n1903) );
  OAI2BB2XL U649 ( .B0(n1573), .B1(n1645), .A0N(\gbuff[27][29] ), .A1N(n1647), 
        .Y(n1902) );
  OAI2BB2XL U650 ( .B0(n1571), .B1(n1645), .A0N(\gbuff[27][30] ), .A1N(n1646), 
        .Y(n1901) );
  OAI2BB2XL U651 ( .B0(n1569), .B1(n1645), .A0N(\gbuff[27][31] ), .A1N(n2800), 
        .Y(n1900) );
  OAI2BB2XL U652 ( .B0(n1585), .B1(n1643), .A0N(\gbuff[28][23] ), .A1N(n1643), 
        .Y(n1876) );
  OAI2BB2XL U653 ( .B0(n1581), .B1(n1643), .A0N(\gbuff[28][25] ), .A1N(n1644), 
        .Y(n1874) );
  OAI2BB2XL U654 ( .B0(n1579), .B1(n1643), .A0N(\gbuff[28][26] ), .A1N(n1644), 
        .Y(n1873) );
  OAI2BB2XL U655 ( .B0(n1577), .B1(n1643), .A0N(\gbuff[28][27] ), .A1N(n1644), 
        .Y(n1872) );
  OAI2BB2XL U656 ( .B0(n1575), .B1(n1643), .A0N(\gbuff[28][28] ), .A1N(n1644), 
        .Y(n1871) );
  OAI2BB2XL U657 ( .B0(n1573), .B1(n1643), .A0N(\gbuff[28][29] ), .A1N(n1644), 
        .Y(n1870) );
  OAI2BB2XL U658 ( .B0(n1571), .B1(n1643), .A0N(\gbuff[28][30] ), .A1N(n1643), 
        .Y(n1869) );
  OAI2BB2XL U659 ( .B0(n1569), .B1(n1643), .A0N(\gbuff[28][31] ), .A1N(n1644), 
        .Y(n1868) );
  OAI2BB2XL U660 ( .B0(n1585), .B1(n1640), .A0N(\gbuff[29][23] ), .A1N(n1640), 
        .Y(n1844) );
  OAI2BB2XL U661 ( .B0(n1581), .B1(n1640), .A0N(\gbuff[29][25] ), .A1N(n1641), 
        .Y(n1842) );
  OAI2BB2XL U662 ( .B0(n1579), .B1(n1640), .A0N(\gbuff[29][26] ), .A1N(n1641), 
        .Y(n1841) );
  OAI2BB2XL U663 ( .B0(n1577), .B1(n1640), .A0N(\gbuff[29][27] ), .A1N(n1641), 
        .Y(n1840) );
  OAI2BB2XL U664 ( .B0(n1575), .B1(n1640), .A0N(\gbuff[29][28] ), .A1N(n1641), 
        .Y(n1839) );
  OAI2BB2XL U665 ( .B0(n1573), .B1(n1640), .A0N(\gbuff[29][29] ), .A1N(n1641), 
        .Y(n1838) );
  OAI2BB2XL U666 ( .B0(n1571), .B1(n1640), .A0N(\gbuff[29][30] ), .A1N(n1640), 
        .Y(n1837) );
  OAI2BB2XL U667 ( .B0(n1569), .B1(n1640), .A0N(\gbuff[29][31] ), .A1N(n1641), 
        .Y(n1836) );
  OAI2BB2XL U668 ( .B0(n1585), .B1(n1637), .A0N(\gbuff[30][23] ), .A1N(n1637), 
        .Y(n1812) );
  OAI2BB2XL U669 ( .B0(n1581), .B1(n1637), .A0N(\gbuff[30][25] ), .A1N(n1638), 
        .Y(n1810) );
  OAI2BB2XL U670 ( .B0(n1579), .B1(n1637), .A0N(\gbuff[30][26] ), .A1N(n1638), 
        .Y(n1809) );
  OAI2BB2XL U671 ( .B0(n1577), .B1(n1637), .A0N(\gbuff[30][27] ), .A1N(n1638), 
        .Y(n1808) );
  OAI2BB2XL U672 ( .B0(n1575), .B1(n1637), .A0N(\gbuff[30][28] ), .A1N(n1638), 
        .Y(n1807) );
  OAI2BB2XL U673 ( .B0(n1573), .B1(n1637), .A0N(\gbuff[30][29] ), .A1N(n1638), 
        .Y(n1806) );
  OAI2BB2XL U674 ( .B0(n1571), .B1(n1637), .A0N(\gbuff[30][30] ), .A1N(n1637), 
        .Y(n1805) );
  OAI2BB2XL U675 ( .B0(n1569), .B1(n1637), .A0N(\gbuff[30][31] ), .A1N(n1638), 
        .Y(n1804) );
  OAI2BB2XL U676 ( .B0(n1585), .B1(n1634), .A0N(\gbuff[31][23] ), .A1N(n1634), 
        .Y(n1780) );
  OAI2BB2XL U677 ( .B0(n1581), .B1(n1634), .A0N(\gbuff[31][25] ), .A1N(n1635), 
        .Y(n1778) );
  OAI2BB2XL U678 ( .B0(n1579), .B1(n1634), .A0N(\gbuff[31][26] ), .A1N(n1635), 
        .Y(n1777) );
  OAI2BB2XL U679 ( .B0(n1577), .B1(n1634), .A0N(\gbuff[31][27] ), .A1N(n1635), 
        .Y(n1776) );
  OAI2BB2XL U680 ( .B0(n1575), .B1(n1634), .A0N(\gbuff[31][28] ), .A1N(n1635), 
        .Y(n1775) );
  OAI2BB2XL U681 ( .B0(n1573), .B1(n1634), .A0N(\gbuff[31][29] ), .A1N(n1635), 
        .Y(n1774) );
  OAI2BB2XL U682 ( .B0(n1571), .B1(n1634), .A0N(\gbuff[31][30] ), .A1N(n1634), 
        .Y(n1773) );
  OAI2BB2XL U683 ( .B0(n1569), .B1(n1634), .A0N(\gbuff[31][31] ), .A1N(n1635), 
        .Y(n1772) );
  OAI2BB2XL U684 ( .B0(n1632), .B1(n1702), .A0N(\gbuff[8][0] ), .A1N(n1703), 
        .Y(n2539) );
  OAI2BB2XL U685 ( .B0(n1630), .B1(n1702), .A0N(\gbuff[8][1] ), .A1N(n10), .Y(
        n2538) );
  OAI2BB2XL U686 ( .B0(n1628), .B1(n1702), .A0N(\gbuff[8][2] ), .A1N(n10), .Y(
        n2537) );
  OAI2BB2XL U687 ( .B0(n1626), .B1(n1702), .A0N(\gbuff[8][3] ), .A1N(n1704), 
        .Y(n2536) );
  OAI2BB2XL U688 ( .B0(n1624), .B1(n1702), .A0N(\gbuff[8][4] ), .A1N(n10), .Y(
        n2535) );
  OAI2BB2XL U689 ( .B0(n1622), .B1(n1702), .A0N(\gbuff[8][5] ), .A1N(n1704), 
        .Y(n2534) );
  OAI2BB2XL U690 ( .B0(n1620), .B1(n1702), .A0N(\gbuff[8][6] ), .A1N(n1704), 
        .Y(n2533) );
  OAI2BB2XL U691 ( .B0(n1618), .B1(n1702), .A0N(\gbuff[8][7] ), .A1N(n1704), 
        .Y(n2532) );
  OAI2BB2XL U692 ( .B0(n1616), .B1(n1702), .A0N(\gbuff[8][8] ), .A1N(n1704), 
        .Y(n2531) );
  OAI2BB2XL U693 ( .B0(n1614), .B1(n1702), .A0N(\gbuff[8][9] ), .A1N(n1704), 
        .Y(n2530) );
  OAI2BB2XL U694 ( .B0(n1612), .B1(n1702), .A0N(\gbuff[8][10] ), .A1N(n1704), 
        .Y(n2529) );
  OAI2BB2XL U695 ( .B0(n1610), .B1(n1702), .A0N(\gbuff[8][11] ), .A1N(n1704), 
        .Y(n2528) );
  OAI2BB2XL U696 ( .B0(n1608), .B1(n1702), .A0N(\gbuff[8][12] ), .A1N(n1704), 
        .Y(n2527) );
  OAI2BB2XL U697 ( .B0(n1606), .B1(n1702), .A0N(\gbuff[8][13] ), .A1N(n1704), 
        .Y(n2526) );
  OAI2BB2XL U698 ( .B0(n1604), .B1(n1702), .A0N(\gbuff[8][14] ), .A1N(n1704), 
        .Y(n2525) );
  OAI2BB2XL U699 ( .B0(n1602), .B1(n1702), .A0N(\gbuff[8][15] ), .A1N(n1703), 
        .Y(n2524) );
  OAI2BB2XL U700 ( .B0(n1600), .B1(n1703), .A0N(\gbuff[8][16] ), .A1N(n1704), 
        .Y(n2523) );
  OAI2BB2XL U701 ( .B0(n1598), .B1(n10), .A0N(\gbuff[8][17] ), .A1N(n1703), 
        .Y(n2522) );
  OAI2BB2XL U702 ( .B0(n1596), .B1(n1702), .A0N(\gbuff[8][18] ), .A1N(n1703), 
        .Y(n2521) );
  OAI2BB2XL U703 ( .B0(n1594), .B1(n1703), .A0N(\gbuff[8][19] ), .A1N(n1703), 
        .Y(n2520) );
  OAI2BB2XL U704 ( .B0(n1592), .B1(n1704), .A0N(\gbuff[8][20] ), .A1N(n1703), 
        .Y(n2519) );
  OAI2BB2XL U705 ( .B0(n1590), .B1(n1703), .A0N(\gbuff[8][21] ), .A1N(n1703), 
        .Y(n2518) );
  OAI2BB2XL U706 ( .B0(n1588), .B1(n1702), .A0N(\gbuff[8][22] ), .A1N(n1704), 
        .Y(n2517) );
  OAI2BB2XL U707 ( .B0(n1584), .B1(n1702), .A0N(\gbuff[8][24] ), .A1N(n1704), 
        .Y(n2515) );
  OAI2BB2XL U708 ( .B0(n1632), .B1(n1699), .A0N(\gbuff[9][0] ), .A1N(n1700), 
        .Y(n2507) );
  OAI2BB2XL U709 ( .B0(n1630), .B1(n1699), .A0N(\gbuff[9][1] ), .A1N(n11), .Y(
        n2506) );
  OAI2BB2XL U710 ( .B0(n1628), .B1(n1699), .A0N(\gbuff[9][2] ), .A1N(n11), .Y(
        n2505) );
  OAI2BB2XL U711 ( .B0(n1626), .B1(n1699), .A0N(\gbuff[9][3] ), .A1N(n1701), 
        .Y(n2504) );
  OAI2BB2XL U712 ( .B0(n1624), .B1(n1699), .A0N(\gbuff[9][4] ), .A1N(n11), .Y(
        n2503) );
  OAI2BB2XL U713 ( .B0(n1622), .B1(n1699), .A0N(\gbuff[9][5] ), .A1N(n1701), 
        .Y(n2502) );
  OAI2BB2XL U714 ( .B0(n1620), .B1(n1699), .A0N(\gbuff[9][6] ), .A1N(n1701), 
        .Y(n2501) );
  OAI2BB2XL U715 ( .B0(n1618), .B1(n1699), .A0N(\gbuff[9][7] ), .A1N(n1701), 
        .Y(n2500) );
  OAI2BB2XL U716 ( .B0(n1616), .B1(n1699), .A0N(\gbuff[9][8] ), .A1N(n1701), 
        .Y(n2499) );
  OAI2BB2XL U717 ( .B0(n1614), .B1(n1699), .A0N(\gbuff[9][9] ), .A1N(n1701), 
        .Y(n2498) );
  OAI2BB2XL U718 ( .B0(n1612), .B1(n1699), .A0N(\gbuff[9][10] ), .A1N(n1701), 
        .Y(n2497) );
  OAI2BB2XL U719 ( .B0(n1610), .B1(n1699), .A0N(\gbuff[9][11] ), .A1N(n1701), 
        .Y(n2496) );
  OAI2BB2XL U720 ( .B0(n1608), .B1(n1699), .A0N(\gbuff[9][12] ), .A1N(n1701), 
        .Y(n2495) );
  OAI2BB2XL U721 ( .B0(n1606), .B1(n1699), .A0N(\gbuff[9][13] ), .A1N(n1701), 
        .Y(n2494) );
  OAI2BB2XL U722 ( .B0(n1604), .B1(n1699), .A0N(\gbuff[9][14] ), .A1N(n1701), 
        .Y(n2493) );
  OAI2BB2XL U723 ( .B0(n1602), .B1(n1699), .A0N(\gbuff[9][15] ), .A1N(n1700), 
        .Y(n2492) );
  OAI2BB2XL U724 ( .B0(n1600), .B1(n1700), .A0N(\gbuff[9][16] ), .A1N(n1701), 
        .Y(n2491) );
  OAI2BB2XL U725 ( .B0(n1598), .B1(n11), .A0N(\gbuff[9][17] ), .A1N(n1700), 
        .Y(n2490) );
  OAI2BB2XL U726 ( .B0(n1596), .B1(n1699), .A0N(\gbuff[9][18] ), .A1N(n1700), 
        .Y(n2489) );
  OAI2BB2XL U727 ( .B0(n1594), .B1(n1700), .A0N(\gbuff[9][19] ), .A1N(n1700), 
        .Y(n2488) );
  OAI2BB2XL U728 ( .B0(n1592), .B1(n1701), .A0N(\gbuff[9][20] ), .A1N(n1700), 
        .Y(n2487) );
  OAI2BB2XL U729 ( .B0(n1590), .B1(n1700), .A0N(\gbuff[9][21] ), .A1N(n1700), 
        .Y(n2486) );
  OAI2BB2XL U730 ( .B0(n1588), .B1(n1699), .A0N(\gbuff[9][22] ), .A1N(n1701), 
        .Y(n2485) );
  OAI2BB2XL U731 ( .B0(n1584), .B1(n1699), .A0N(\gbuff[9][24] ), .A1N(n1701), 
        .Y(n2483) );
  OAI2BB2XL U732 ( .B0(n1632), .B1(n1697), .A0N(\gbuff[10][0] ), .A1N(n1696), 
        .Y(n2475) );
  OAI2BB2XL U733 ( .B0(n1630), .B1(n1696), .A0N(\gbuff[10][1] ), .A1N(n1697), 
        .Y(n2474) );
  OAI2BB2XL U734 ( .B0(n1628), .B1(n1696), .A0N(\gbuff[10][2] ), .A1N(n1696), 
        .Y(n2473) );
  OAI2BB2XL U735 ( .B0(n1626), .B1(n1696), .A0N(\gbuff[10][3] ), .A1N(n1698), 
        .Y(n2472) );
  OAI2BB2XL U736 ( .B0(n1624), .B1(n1696), .A0N(\gbuff[10][4] ), .A1N(n1697), 
        .Y(n2471) );
  OAI2BB2XL U737 ( .B0(n1622), .B1(n1696), .A0N(\gbuff[10][5] ), .A1N(n1698), 
        .Y(n2470) );
  OAI2BB2XL U738 ( .B0(n1620), .B1(n1696), .A0N(\gbuff[10][6] ), .A1N(n1698), 
        .Y(n2469) );
  OAI2BB2XL U739 ( .B0(n1618), .B1(n1696), .A0N(\gbuff[10][7] ), .A1N(n1698), 
        .Y(n2468) );
  OAI2BB2XL U740 ( .B0(n1616), .B1(n1696), .A0N(\gbuff[10][8] ), .A1N(n1698), 
        .Y(n2467) );
  OAI2BB2XL U741 ( .B0(n1614), .B1(n1696), .A0N(\gbuff[10][9] ), .A1N(n1698), 
        .Y(n2466) );
  OAI2BB2XL U742 ( .B0(n1612), .B1(n1696), .A0N(\gbuff[10][10] ), .A1N(n1698), 
        .Y(n2465) );
  OAI2BB2XL U743 ( .B0(n1610), .B1(n1696), .A0N(\gbuff[10][11] ), .A1N(n1698), 
        .Y(n2464) );
  OAI2BB2XL U744 ( .B0(n1608), .B1(n1696), .A0N(\gbuff[10][12] ), .A1N(n1698), 
        .Y(n2463) );
  OAI2BB2XL U745 ( .B0(n1606), .B1(n1697), .A0N(\gbuff[10][13] ), .A1N(n1698), 
        .Y(n2462) );
  OAI2BB2XL U746 ( .B0(n1604), .B1(n1697), .A0N(\gbuff[10][14] ), .A1N(n1698), 
        .Y(n2461) );
  OAI2BB2XL U747 ( .B0(n1602), .B1(n1697), .A0N(\gbuff[10][15] ), .A1N(n1698), 
        .Y(n2460) );
  OAI2BB2XL U748 ( .B0(n1600), .B1(n1697), .A0N(\gbuff[10][16] ), .A1N(n1698), 
        .Y(n2459) );
  OAI2BB2XL U749 ( .B0(n1598), .B1(n1697), .A0N(\gbuff[10][17] ), .A1N(n13), 
        .Y(n2458) );
  OAI2BB2XL U750 ( .B0(n1596), .B1(n1697), .A0N(\gbuff[10][18] ), .A1N(n13), 
        .Y(n2457) );
  OAI2BB2XL U751 ( .B0(n1594), .B1(n1697), .A0N(\gbuff[10][19] ), .A1N(n1698), 
        .Y(n2456) );
  OAI2BB2XL U752 ( .B0(n1592), .B1(n1697), .A0N(\gbuff[10][20] ), .A1N(n1698), 
        .Y(n2455) );
  OAI2BB2XL U753 ( .B0(n1590), .B1(n1697), .A0N(\gbuff[10][21] ), .A1N(n1696), 
        .Y(n2454) );
  OAI2BB2XL U754 ( .B0(n1588), .B1(n1697), .A0N(\gbuff[10][22] ), .A1N(n1698), 
        .Y(n2453) );
  OAI2BB2XL U755 ( .B0(n1584), .B1(n1697), .A0N(\gbuff[10][24] ), .A1N(n1698), 
        .Y(n2451) );
  OAI2BB2XL U756 ( .B0(n1632), .B1(n1693), .A0N(\gbuff[11][0] ), .A1N(n1693), 
        .Y(n2443) );
  OAI2BB2XL U757 ( .B0(n1630), .B1(n1694), .A0N(\gbuff[11][1] ), .A1N(n1693), 
        .Y(n2442) );
  OAI2BB2XL U758 ( .B0(n1628), .B1(n1694), .A0N(\gbuff[11][2] ), .A1N(n1693), 
        .Y(n2441) );
  OAI2BB2XL U759 ( .B0(n1626), .B1(n1694), .A0N(\gbuff[11][3] ), .A1N(n1695), 
        .Y(n2440) );
  OAI2BB2XL U760 ( .B0(n1624), .B1(n1694), .A0N(\gbuff[11][4] ), .A1N(n1693), 
        .Y(n2439) );
  OAI2BB2XL U761 ( .B0(n1622), .B1(n1694), .A0N(\gbuff[11][5] ), .A1N(n1695), 
        .Y(n2438) );
  OAI2BB2XL U762 ( .B0(n1620), .B1(n1694), .A0N(\gbuff[11][6] ), .A1N(n1695), 
        .Y(n2437) );
  OAI2BB2XL U763 ( .B0(n1618), .B1(n1694), .A0N(\gbuff[11][7] ), .A1N(n1695), 
        .Y(n2436) );
  OAI2BB2XL U764 ( .B0(n1616), .B1(n1694), .A0N(\gbuff[11][8] ), .A1N(n1695), 
        .Y(n2435) );
  OAI2BB2XL U765 ( .B0(n1614), .B1(n1694), .A0N(\gbuff[11][9] ), .A1N(n1695), 
        .Y(n2434) );
  OAI2BB2XL U766 ( .B0(n1612), .B1(n1694), .A0N(\gbuff[11][10] ), .A1N(n1695), 
        .Y(n2433) );
  OAI2BB2XL U767 ( .B0(n1610), .B1(n1694), .A0N(\gbuff[11][11] ), .A1N(n1695), 
        .Y(n2432) );
  OAI2BB2XL U768 ( .B0(n1608), .B1(n1694), .A0N(\gbuff[11][12] ), .A1N(n1695), 
        .Y(n2431) );
  OAI2BB2XL U769 ( .B0(n1606), .B1(n1693), .A0N(\gbuff[11][13] ), .A1N(n1695), 
        .Y(n2430) );
  OAI2BB2XL U770 ( .B0(n1604), .B1(n1693), .A0N(\gbuff[11][14] ), .A1N(n1695), 
        .Y(n2429) );
  OAI2BB2XL U771 ( .B0(n1602), .B1(n1693), .A0N(\gbuff[11][15] ), .A1N(n6), 
        .Y(n2428) );
  OAI2BB2XL U772 ( .B0(n1600), .B1(n1693), .A0N(\gbuff[11][16] ), .A1N(n1695), 
        .Y(n2427) );
  OAI2BB2XL U773 ( .B0(n1598), .B1(n1693), .A0N(\gbuff[11][17] ), .A1N(n1693), 
        .Y(n2426) );
  OAI2BB2XL U774 ( .B0(n1596), .B1(n1693), .A0N(\gbuff[11][18] ), .A1N(n1693), 
        .Y(n2425) );
  OAI2BB2XL U775 ( .B0(n1594), .B1(n1693), .A0N(\gbuff[11][19] ), .A1N(n1693), 
        .Y(n2424) );
  OAI2BB2XL U776 ( .B0(n1592), .B1(n1693), .A0N(\gbuff[11][20] ), .A1N(n1693), 
        .Y(n2423) );
  OAI2BB2XL U777 ( .B0(n1590), .B1(n1694), .A0N(\gbuff[11][21] ), .A1N(n1693), 
        .Y(n2422) );
  OAI2BB2XL U778 ( .B0(n1588), .B1(n1693), .A0N(\gbuff[11][22] ), .A1N(n1695), 
        .Y(n2421) );
  OAI2BB2XL U779 ( .B0(n1584), .B1(n1694), .A0N(\gbuff[11][24] ), .A1N(n1695), 
        .Y(n2419) );
  OAI2BB2XL U780 ( .B0(n1632), .B1(n1690), .A0N(\gbuff[12][0] ), .A1N(n1691), 
        .Y(n2411) );
  OAI2BB2XL U781 ( .B0(n1630), .B1(n1690), .A0N(\gbuff[12][1] ), .A1N(n12), 
        .Y(n2410) );
  OAI2BB2XL U782 ( .B0(n1628), .B1(n1690), .A0N(\gbuff[12][2] ), .A1N(n12), 
        .Y(n2409) );
  OAI2BB2XL U783 ( .B0(n1626), .B1(n1690), .A0N(\gbuff[12][3] ), .A1N(n1692), 
        .Y(n2408) );
  OAI2BB2XL U784 ( .B0(n1624), .B1(n1690), .A0N(\gbuff[12][4] ), .A1N(n12), 
        .Y(n2407) );
  OAI2BB2XL U785 ( .B0(n1622), .B1(n1690), .A0N(\gbuff[12][5] ), .A1N(n1692), 
        .Y(n2406) );
  OAI2BB2XL U786 ( .B0(n1620), .B1(n1690), .A0N(\gbuff[12][6] ), .A1N(n1692), 
        .Y(n2405) );
  OAI2BB2XL U787 ( .B0(n1618), .B1(n1690), .A0N(\gbuff[12][7] ), .A1N(n1692), 
        .Y(n2404) );
  OAI2BB2XL U788 ( .B0(n1616), .B1(n1690), .A0N(\gbuff[12][8] ), .A1N(n1692), 
        .Y(n2403) );
  OAI2BB2XL U789 ( .B0(n1614), .B1(n1690), .A0N(\gbuff[12][9] ), .A1N(n1692), 
        .Y(n2402) );
  OAI2BB2XL U790 ( .B0(n1612), .B1(n1690), .A0N(\gbuff[12][10] ), .A1N(n1692), 
        .Y(n2401) );
  OAI2BB2XL U791 ( .B0(n1610), .B1(n1690), .A0N(\gbuff[12][11] ), .A1N(n1692), 
        .Y(n2400) );
  OAI2BB2XL U792 ( .B0(n1608), .B1(n1690), .A0N(\gbuff[12][12] ), .A1N(n1692), 
        .Y(n2399) );
  OAI2BB2XL U793 ( .B0(n1606), .B1(n1690), .A0N(\gbuff[12][13] ), .A1N(n1692), 
        .Y(n2398) );
  OAI2BB2XL U794 ( .B0(n1604), .B1(n1690), .A0N(\gbuff[12][14] ), .A1N(n1692), 
        .Y(n2397) );
  OAI2BB2XL U795 ( .B0(n1602), .B1(n1690), .A0N(\gbuff[12][15] ), .A1N(n1691), 
        .Y(n2396) );
  OAI2BB2XL U796 ( .B0(n1600), .B1(n1691), .A0N(\gbuff[12][16] ), .A1N(n1692), 
        .Y(n2395) );
  OAI2BB2XL U797 ( .B0(n1598), .B1(n12), .A0N(\gbuff[12][17] ), .A1N(n1691), 
        .Y(n2394) );
  OAI2BB2XL U798 ( .B0(n1596), .B1(n1690), .A0N(\gbuff[12][18] ), .A1N(n1691), 
        .Y(n2393) );
  OAI2BB2XL U799 ( .B0(n1594), .B1(n1691), .A0N(\gbuff[12][19] ), .A1N(n1691), 
        .Y(n2392) );
  OAI2BB2XL U800 ( .B0(n1592), .B1(n1692), .A0N(\gbuff[12][20] ), .A1N(n1691), 
        .Y(n2391) );
  OAI2BB2XL U801 ( .B0(n1590), .B1(n1691), .A0N(\gbuff[12][21] ), .A1N(n1691), 
        .Y(n2390) );
  OAI2BB2XL U802 ( .B0(n1588), .B1(n1690), .A0N(\gbuff[12][22] ), .A1N(n1692), 
        .Y(n2389) );
  OAI2BB2XL U803 ( .B0(n1584), .B1(n1690), .A0N(\gbuff[12][24] ), .A1N(n1692), 
        .Y(n2387) );
  OAI2BB2XL U804 ( .B0(n1632), .B1(n1687), .A0N(\gbuff[13][0] ), .A1N(n1687), 
        .Y(n2379) );
  OAI2BB2XL U805 ( .B0(n1630), .B1(n1688), .A0N(\gbuff[13][1] ), .A1N(n1687), 
        .Y(n2378) );
  OAI2BB2XL U806 ( .B0(n1628), .B1(n1688), .A0N(\gbuff[13][2] ), .A1N(n1687), 
        .Y(n2377) );
  OAI2BB2XL U807 ( .B0(n1626), .B1(n1688), .A0N(\gbuff[13][3] ), .A1N(n1689), 
        .Y(n2376) );
  OAI2BB2XL U808 ( .B0(n1624), .B1(n1688), .A0N(\gbuff[13][4] ), .A1N(n1687), 
        .Y(n2375) );
  OAI2BB2XL U809 ( .B0(n1622), .B1(n1688), .A0N(\gbuff[13][5] ), .A1N(n1689), 
        .Y(n2374) );
  OAI2BB2XL U810 ( .B0(n1620), .B1(n1688), .A0N(\gbuff[13][6] ), .A1N(n1689), 
        .Y(n2373) );
  OAI2BB2XL U811 ( .B0(n1618), .B1(n1688), .A0N(\gbuff[13][7] ), .A1N(n1689), 
        .Y(n2372) );
  OAI2BB2XL U812 ( .B0(n1616), .B1(n1688), .A0N(\gbuff[13][8] ), .A1N(n1689), 
        .Y(n2371) );
  OAI2BB2XL U813 ( .B0(n1614), .B1(n1688), .A0N(\gbuff[13][9] ), .A1N(n1689), 
        .Y(n2370) );
  OAI2BB2XL U814 ( .B0(n1612), .B1(n1688), .A0N(\gbuff[13][10] ), .A1N(n1689), 
        .Y(n2369) );
  OAI2BB2XL U815 ( .B0(n1610), .B1(n1688), .A0N(\gbuff[13][11] ), .A1N(n1689), 
        .Y(n2368) );
  OAI2BB2XL U816 ( .B0(n1608), .B1(n1688), .A0N(\gbuff[13][12] ), .A1N(n1689), 
        .Y(n2367) );
  OAI2BB2XL U817 ( .B0(n1606), .B1(n1687), .A0N(\gbuff[13][13] ), .A1N(n1689), 
        .Y(n2366) );
  OAI2BB2XL U818 ( .B0(n1604), .B1(n1687), .A0N(\gbuff[13][14] ), .A1N(n1689), 
        .Y(n2365) );
  OAI2BB2XL U819 ( .B0(n1602), .B1(n1687), .A0N(\gbuff[13][15] ), .A1N(n7), 
        .Y(n2364) );
  OAI2BB2XL U820 ( .B0(n1600), .B1(n1687), .A0N(\gbuff[13][16] ), .A1N(n1689), 
        .Y(n2363) );
  OAI2BB2XL U821 ( .B0(n1598), .B1(n1687), .A0N(\gbuff[13][17] ), .A1N(n1687), 
        .Y(n2362) );
  OAI2BB2XL U822 ( .B0(n1596), .B1(n1687), .A0N(\gbuff[13][18] ), .A1N(n1687), 
        .Y(n2361) );
  OAI2BB2XL U823 ( .B0(n1594), .B1(n1687), .A0N(\gbuff[13][19] ), .A1N(n1687), 
        .Y(n2360) );
  OAI2BB2XL U824 ( .B0(n1592), .B1(n1687), .A0N(\gbuff[13][20] ), .A1N(n1687), 
        .Y(n2359) );
  OAI2BB2XL U825 ( .B0(n1590), .B1(n1688), .A0N(\gbuff[13][21] ), .A1N(n1687), 
        .Y(n2358) );
  OAI2BB2XL U826 ( .B0(n1588), .B1(n1687), .A0N(\gbuff[13][22] ), .A1N(n1689), 
        .Y(n2357) );
  OAI2BB2XL U827 ( .B0(n1584), .B1(n1688), .A0N(\gbuff[13][24] ), .A1N(n1689), 
        .Y(n2355) );
  OAI2BB2XL U828 ( .B0(n1632), .B1(n1684), .A0N(\gbuff[14][0] ), .A1N(n1684), 
        .Y(n2347) );
  OAI2BB2XL U829 ( .B0(n1630), .B1(n1685), .A0N(\gbuff[14][1] ), .A1N(n1684), 
        .Y(n2346) );
  OAI2BB2XL U830 ( .B0(n1628), .B1(n1685), .A0N(\gbuff[14][2] ), .A1N(n1684), 
        .Y(n2345) );
  OAI2BB2XL U831 ( .B0(n1626), .B1(n1685), .A0N(\gbuff[14][3] ), .A1N(n1686), 
        .Y(n2344) );
  OAI2BB2XL U832 ( .B0(n1624), .B1(n1685), .A0N(\gbuff[14][4] ), .A1N(n1684), 
        .Y(n2343) );
  OAI2BB2XL U833 ( .B0(n1622), .B1(n1685), .A0N(\gbuff[14][5] ), .A1N(n1686), 
        .Y(n2342) );
  OAI2BB2XL U834 ( .B0(n1620), .B1(n1685), .A0N(\gbuff[14][6] ), .A1N(n1686), 
        .Y(n2341) );
  OAI2BB2XL U835 ( .B0(n1618), .B1(n1685), .A0N(\gbuff[14][7] ), .A1N(n1686), 
        .Y(n2340) );
  OAI2BB2XL U836 ( .B0(n1616), .B1(n1685), .A0N(\gbuff[14][8] ), .A1N(n1686), 
        .Y(n2339) );
  OAI2BB2XL U837 ( .B0(n1614), .B1(n1685), .A0N(\gbuff[14][9] ), .A1N(n1686), 
        .Y(n2338) );
  OAI2BB2XL U838 ( .B0(n1612), .B1(n1685), .A0N(\gbuff[14][10] ), .A1N(n1686), 
        .Y(n2337) );
  OAI2BB2XL U839 ( .B0(n1610), .B1(n1685), .A0N(\gbuff[14][11] ), .A1N(n1686), 
        .Y(n2336) );
  OAI2BB2XL U840 ( .B0(n1608), .B1(n1685), .A0N(\gbuff[14][12] ), .A1N(n1686), 
        .Y(n2335) );
  OAI2BB2XL U841 ( .B0(n1606), .B1(n1684), .A0N(\gbuff[14][13] ), .A1N(n1686), 
        .Y(n2334) );
  OAI2BB2XL U842 ( .B0(n1604), .B1(n1684), .A0N(\gbuff[14][14] ), .A1N(n1686), 
        .Y(n2333) );
  OAI2BB2XL U843 ( .B0(n1602), .B1(n1684), .A0N(\gbuff[14][15] ), .A1N(n8), 
        .Y(n2332) );
  OAI2BB2XL U844 ( .B0(n1600), .B1(n1684), .A0N(\gbuff[14][16] ), .A1N(n1686), 
        .Y(n2331) );
  OAI2BB2XL U845 ( .B0(n1598), .B1(n1684), .A0N(\gbuff[14][17] ), .A1N(n1684), 
        .Y(n2330) );
  OAI2BB2XL U846 ( .B0(n1596), .B1(n1684), .A0N(\gbuff[14][18] ), .A1N(n1684), 
        .Y(n2329) );
  OAI2BB2XL U847 ( .B0(n1594), .B1(n1684), .A0N(\gbuff[14][19] ), .A1N(n1684), 
        .Y(n2328) );
  OAI2BB2XL U848 ( .B0(n1592), .B1(n1684), .A0N(\gbuff[14][20] ), .A1N(n1684), 
        .Y(n2327) );
  OAI2BB2XL U849 ( .B0(n1590), .B1(n1685), .A0N(\gbuff[14][21] ), .A1N(n1684), 
        .Y(n2326) );
  OAI2BB2XL U850 ( .B0(n1588), .B1(n1684), .A0N(\gbuff[14][22] ), .A1N(n1686), 
        .Y(n2325) );
  OAI2BB2XL U851 ( .B0(n1584), .B1(n1685), .A0N(\gbuff[14][24] ), .A1N(n1686), 
        .Y(n2323) );
  OAI2BB2XL U852 ( .B0(n1632), .B1(n1681), .A0N(\gbuff[15][0] ), .A1N(n1681), 
        .Y(n2315) );
  OAI2BB2XL U853 ( .B0(n1630), .B1(n1682), .A0N(\gbuff[15][1] ), .A1N(n1681), 
        .Y(n2314) );
  OAI2BB2XL U854 ( .B0(n1628), .B1(n1682), .A0N(\gbuff[15][2] ), .A1N(n1681), 
        .Y(n2313) );
  OAI2BB2XL U855 ( .B0(n1626), .B1(n1682), .A0N(\gbuff[15][3] ), .A1N(n1683), 
        .Y(n2312) );
  OAI2BB2XL U856 ( .B0(n1624), .B1(n1682), .A0N(\gbuff[15][4] ), .A1N(n1681), 
        .Y(n2311) );
  OAI2BB2XL U857 ( .B0(n1622), .B1(n1682), .A0N(\gbuff[15][5] ), .A1N(n1683), 
        .Y(n2310) );
  OAI2BB2XL U858 ( .B0(n1620), .B1(n1682), .A0N(\gbuff[15][6] ), .A1N(n1683), 
        .Y(n2309) );
  OAI2BB2XL U859 ( .B0(n1618), .B1(n1682), .A0N(\gbuff[15][7] ), .A1N(n1683), 
        .Y(n2308) );
  OAI2BB2XL U860 ( .B0(n1616), .B1(n1682), .A0N(\gbuff[15][8] ), .A1N(n1683), 
        .Y(n2307) );
  OAI2BB2XL U861 ( .B0(n1614), .B1(n1682), .A0N(\gbuff[15][9] ), .A1N(n1683), 
        .Y(n2306) );
  OAI2BB2XL U862 ( .B0(n1612), .B1(n1682), .A0N(\gbuff[15][10] ), .A1N(n1683), 
        .Y(n2305) );
  OAI2BB2XL U863 ( .B0(n1610), .B1(n1682), .A0N(\gbuff[15][11] ), .A1N(n1683), 
        .Y(n2304) );
  OAI2BB2XL U864 ( .B0(n1608), .B1(n1682), .A0N(\gbuff[15][12] ), .A1N(n1683), 
        .Y(n2303) );
  OAI2BB2XL U865 ( .B0(n1606), .B1(n1681), .A0N(\gbuff[15][13] ), .A1N(n1683), 
        .Y(n2302) );
  OAI2BB2XL U866 ( .B0(n1604), .B1(n1681), .A0N(\gbuff[15][14] ), .A1N(n1683), 
        .Y(n2301) );
  OAI2BB2XL U867 ( .B0(n1602), .B1(n1681), .A0N(\gbuff[15][15] ), .A1N(n9), 
        .Y(n2300) );
  OAI2BB2XL U868 ( .B0(n1600), .B1(n1681), .A0N(\gbuff[15][16] ), .A1N(n1683), 
        .Y(n2299) );
  OAI2BB2XL U869 ( .B0(n1598), .B1(n1681), .A0N(\gbuff[15][17] ), .A1N(n1681), 
        .Y(n2298) );
  OAI2BB2XL U870 ( .B0(n1596), .B1(n1681), .A0N(\gbuff[15][18] ), .A1N(n1681), 
        .Y(n2297) );
  OAI2BB2XL U871 ( .B0(n1594), .B1(n1681), .A0N(\gbuff[15][19] ), .A1N(n1681), 
        .Y(n2296) );
  OAI2BB2XL U872 ( .B0(n1592), .B1(n1681), .A0N(\gbuff[15][20] ), .A1N(n1681), 
        .Y(n2295) );
  OAI2BB2XL U873 ( .B0(n1590), .B1(n1682), .A0N(\gbuff[15][21] ), .A1N(n1681), 
        .Y(n2294) );
  OAI2BB2XL U874 ( .B0(n1588), .B1(n1681), .A0N(\gbuff[15][22] ), .A1N(n1683), 
        .Y(n2293) );
  OAI2BB2XL U875 ( .B0(n1584), .B1(n1682), .A0N(\gbuff[15][24] ), .A1N(n1683), 
        .Y(n2291) );
  OAI2BB2XL U876 ( .B0(n1632), .B1(n1679), .A0N(\gbuff[16][0] ), .A1N(n1678), 
        .Y(n2283) );
  OAI2BB2XL U877 ( .B0(n1630), .B1(n1679), .A0N(\gbuff[16][1] ), .A1N(n1678), 
        .Y(n2282) );
  OAI2BB2XL U878 ( .B0(n1628), .B1(n1679), .A0N(\gbuff[16][2] ), .A1N(n1678), 
        .Y(n2281) );
  OAI2BB2XL U879 ( .B0(n1626), .B1(n1679), .A0N(\gbuff[16][3] ), .A1N(n1680), 
        .Y(n2280) );
  OAI2BB2XL U880 ( .B0(n1624), .B1(n1679), .A0N(\gbuff[16][4] ), .A1N(n1678), 
        .Y(n2279) );
  OAI2BB2XL U881 ( .B0(n1622), .B1(n1679), .A0N(\gbuff[16][5] ), .A1N(n1680), 
        .Y(n2278) );
  OAI2BB2XL U882 ( .B0(n1620), .B1(n1679), .A0N(\gbuff[16][6] ), .A1N(n1680), 
        .Y(n2277) );
  OAI2BB2XL U883 ( .B0(n1618), .B1(n1679), .A0N(\gbuff[16][7] ), .A1N(n1680), 
        .Y(n2276) );
  OAI2BB2XL U884 ( .B0(n1616), .B1(n1679), .A0N(\gbuff[16][8] ), .A1N(n1680), 
        .Y(n2275) );
  OAI2BB2XL U885 ( .B0(n1614), .B1(n1679), .A0N(\gbuff[16][9] ), .A1N(n1680), 
        .Y(n2274) );
  OAI2BB2XL U886 ( .B0(n1612), .B1(n1679), .A0N(\gbuff[16][10] ), .A1N(n1680), 
        .Y(n2273) );
  OAI2BB2XL U887 ( .B0(n1610), .B1(n1679), .A0N(\gbuff[16][11] ), .A1N(n1680), 
        .Y(n2272) );
  OAI2BB2XL U888 ( .B0(n1608), .B1(n1679), .A0N(\gbuff[16][12] ), .A1N(n1680), 
        .Y(n2271) );
  OAI2BB2XL U889 ( .B0(n1606), .B1(n1679), .A0N(\gbuff[16][13] ), .A1N(n1680), 
        .Y(n2270) );
  OAI2BB2XL U890 ( .B0(n1604), .B1(n1679), .A0N(\gbuff[16][14] ), .A1N(n1680), 
        .Y(n2269) );
  OAI2BB2XL U891 ( .B0(n1602), .B1(n1679), .A0N(\gbuff[16][15] ), .A1N(n1678), 
        .Y(n2268) );
  OAI2BB2XL U892 ( .B0(n1600), .B1(n1678), .A0N(\gbuff[16][16] ), .A1N(n1680), 
        .Y(n2267) );
  OAI2BB2XL U893 ( .B0(n1598), .B1(n1678), .A0N(\gbuff[16][17] ), .A1N(n1680), 
        .Y(n2266) );
  OAI2BB2XL U894 ( .B0(n1596), .B1(n2813), .A0N(\gbuff[16][18] ), .A1N(n1678), 
        .Y(n2265) );
  OAI2BB2XL U895 ( .B0(n1594), .B1(n1679), .A0N(\gbuff[16][19] ), .A1N(n1678), 
        .Y(n2264) );
  OAI2BB2XL U896 ( .B0(n1592), .B1(n2813), .A0N(\gbuff[16][20] ), .A1N(n1678), 
        .Y(n2263) );
  OAI2BB2XL U897 ( .B0(n1590), .B1(n2813), .A0N(\gbuff[16][21] ), .A1N(n1678), 
        .Y(n2262) );
  OAI2BB2XL U898 ( .B0(n1588), .B1(n1678), .A0N(\gbuff[16][22] ), .A1N(n1680), 
        .Y(n2261) );
  OAI2BB2XL U899 ( .B0(n1584), .B1(n2813), .A0N(\gbuff[16][24] ), .A1N(n1680), 
        .Y(n2259) );
  OAI2BB2XL U900 ( .B0(n1632), .B1(n1676), .A0N(\gbuff[17][0] ), .A1N(n1675), 
        .Y(n2251) );
  OAI2BB2XL U901 ( .B0(n1630), .B1(n1676), .A0N(\gbuff[17][1] ), .A1N(n1675), 
        .Y(n2250) );
  OAI2BB2XL U902 ( .B0(n1628), .B1(n1676), .A0N(\gbuff[17][2] ), .A1N(n1675), 
        .Y(n2249) );
  OAI2BB2XL U903 ( .B0(n1626), .B1(n1676), .A0N(\gbuff[17][3] ), .A1N(n1677), 
        .Y(n2248) );
  OAI2BB2XL U904 ( .B0(n1624), .B1(n1676), .A0N(\gbuff[17][4] ), .A1N(n1675), 
        .Y(n2247) );
  OAI2BB2XL U905 ( .B0(n1622), .B1(n1676), .A0N(\gbuff[17][5] ), .A1N(n1677), 
        .Y(n2246) );
  OAI2BB2XL U906 ( .B0(n1620), .B1(n1676), .A0N(\gbuff[17][6] ), .A1N(n1677), 
        .Y(n2245) );
  OAI2BB2XL U907 ( .B0(n1618), .B1(n1676), .A0N(\gbuff[17][7] ), .A1N(n1677), 
        .Y(n2244) );
  OAI2BB2XL U908 ( .B0(n1616), .B1(n1676), .A0N(\gbuff[17][8] ), .A1N(n1677), 
        .Y(n2243) );
  OAI2BB2XL U909 ( .B0(n1614), .B1(n1676), .A0N(\gbuff[17][9] ), .A1N(n1677), 
        .Y(n2242) );
  OAI2BB2XL U910 ( .B0(n1612), .B1(n1676), .A0N(\gbuff[17][10] ), .A1N(n1677), 
        .Y(n2241) );
  OAI2BB2XL U911 ( .B0(n1610), .B1(n1676), .A0N(\gbuff[17][11] ), .A1N(n1677), 
        .Y(n2240) );
  OAI2BB2XL U912 ( .B0(n1608), .B1(n1676), .A0N(\gbuff[17][12] ), .A1N(n1677), 
        .Y(n2239) );
  OAI2BB2XL U913 ( .B0(n1606), .B1(n1676), .A0N(\gbuff[17][13] ), .A1N(n1677), 
        .Y(n2238) );
  OAI2BB2XL U914 ( .B0(n1604), .B1(n1676), .A0N(\gbuff[17][14] ), .A1N(n1677), 
        .Y(n2237) );
  OAI2BB2XL U915 ( .B0(n1602), .B1(n1676), .A0N(\gbuff[17][15] ), .A1N(n1675), 
        .Y(n2236) );
  OAI2BB2XL U916 ( .B0(n1600), .B1(n1675), .A0N(\gbuff[17][16] ), .A1N(n1677), 
        .Y(n2235) );
  OAI2BB2XL U917 ( .B0(n1598), .B1(n1675), .A0N(\gbuff[17][17] ), .A1N(n1677), 
        .Y(n2234) );
  OAI2BB2XL U918 ( .B0(n1596), .B1(n2811), .A0N(\gbuff[17][18] ), .A1N(n1675), 
        .Y(n2233) );
  OAI2BB2XL U919 ( .B0(n1594), .B1(n1676), .A0N(\gbuff[17][19] ), .A1N(n1675), 
        .Y(n2232) );
  OAI2BB2XL U920 ( .B0(n1592), .B1(n2811), .A0N(\gbuff[17][20] ), .A1N(n1675), 
        .Y(n2231) );
  OAI2BB2XL U921 ( .B0(n1590), .B1(n2811), .A0N(\gbuff[17][21] ), .A1N(n1675), 
        .Y(n2230) );
  OAI2BB2XL U922 ( .B0(n1588), .B1(n1675), .A0N(\gbuff[17][22] ), .A1N(n1677), 
        .Y(n2229) );
  OAI2BB2XL U923 ( .B0(n1584), .B1(n2811), .A0N(\gbuff[17][24] ), .A1N(n1677), 
        .Y(n2227) );
  OAI2BB2XL U924 ( .B0(n1632), .B1(n1673), .A0N(\gbuff[18][0] ), .A1N(n1672), 
        .Y(n2219) );
  OAI2BB2XL U925 ( .B0(n1630), .B1(n1673), .A0N(\gbuff[18][1] ), .A1N(n1672), 
        .Y(n2218) );
  OAI2BB2XL U926 ( .B0(n1628), .B1(n1673), .A0N(\gbuff[18][2] ), .A1N(n1672), 
        .Y(n2217) );
  OAI2BB2XL U927 ( .B0(n1626), .B1(n1673), .A0N(\gbuff[18][3] ), .A1N(n1674), 
        .Y(n2216) );
  OAI2BB2XL U928 ( .B0(n1624), .B1(n1673), .A0N(\gbuff[18][4] ), .A1N(n1672), 
        .Y(n2215) );
  OAI2BB2XL U929 ( .B0(n1622), .B1(n1673), .A0N(\gbuff[18][5] ), .A1N(n1674), 
        .Y(n2214) );
  OAI2BB2XL U930 ( .B0(n1620), .B1(n1673), .A0N(\gbuff[18][6] ), .A1N(n1674), 
        .Y(n2213) );
  OAI2BB2XL U931 ( .B0(n1618), .B1(n1673), .A0N(\gbuff[18][7] ), .A1N(n1674), 
        .Y(n2212) );
  OAI2BB2XL U932 ( .B0(n1616), .B1(n1673), .A0N(\gbuff[18][8] ), .A1N(n1674), 
        .Y(n2211) );
  OAI2BB2XL U933 ( .B0(n1614), .B1(n1673), .A0N(\gbuff[18][9] ), .A1N(n1674), 
        .Y(n2210) );
  OAI2BB2XL U934 ( .B0(n1612), .B1(n1673), .A0N(\gbuff[18][10] ), .A1N(n1674), 
        .Y(n2209) );
  OAI2BB2XL U935 ( .B0(n1610), .B1(n1673), .A0N(\gbuff[18][11] ), .A1N(n1674), 
        .Y(n2208) );
  OAI2BB2XL U936 ( .B0(n1608), .B1(n1673), .A0N(\gbuff[18][12] ), .A1N(n1674), 
        .Y(n2207) );
  OAI2BB2XL U937 ( .B0(n1606), .B1(n1673), .A0N(\gbuff[18][13] ), .A1N(n1674), 
        .Y(n2206) );
  OAI2BB2XL U938 ( .B0(n1604), .B1(n1673), .A0N(\gbuff[18][14] ), .A1N(n1674), 
        .Y(n2205) );
  OAI2BB2XL U939 ( .B0(n1602), .B1(n1673), .A0N(\gbuff[18][15] ), .A1N(n1672), 
        .Y(n2204) );
  OAI2BB2XL U940 ( .B0(n1600), .B1(n1672), .A0N(\gbuff[18][16] ), .A1N(n1674), 
        .Y(n2203) );
  OAI2BB2XL U941 ( .B0(n1598), .B1(n1672), .A0N(\gbuff[18][17] ), .A1N(n1674), 
        .Y(n2202) );
  OAI2BB2XL U942 ( .B0(n1596), .B1(n2810), .A0N(\gbuff[18][18] ), .A1N(n1672), 
        .Y(n2201) );
  OAI2BB2XL U943 ( .B0(n1594), .B1(n1673), .A0N(\gbuff[18][19] ), .A1N(n1672), 
        .Y(n2200) );
  OAI2BB2XL U944 ( .B0(n1592), .B1(n2810), .A0N(\gbuff[18][20] ), .A1N(n1672), 
        .Y(n2199) );
  OAI2BB2XL U945 ( .B0(n1590), .B1(n2810), .A0N(\gbuff[18][21] ), .A1N(n1672), 
        .Y(n2198) );
  OAI2BB2XL U946 ( .B0(n1588), .B1(n1672), .A0N(\gbuff[18][22] ), .A1N(n1674), 
        .Y(n2197) );
  OAI2BB2XL U947 ( .B0(n1584), .B1(n2810), .A0N(\gbuff[18][24] ), .A1N(n1674), 
        .Y(n2195) );
  OAI2BB2XL U948 ( .B0(n1632), .B1(n1670), .A0N(\gbuff[19][0] ), .A1N(n1669), 
        .Y(n2187) );
  OAI2BB2XL U949 ( .B0(n1630), .B1(n1670), .A0N(\gbuff[19][1] ), .A1N(n1669), 
        .Y(n2186) );
  OAI2BB2XL U950 ( .B0(n1628), .B1(n1670), .A0N(\gbuff[19][2] ), .A1N(n1669), 
        .Y(n2185) );
  OAI2BB2XL U951 ( .B0(n1626), .B1(n1670), .A0N(\gbuff[19][3] ), .A1N(n1671), 
        .Y(n2184) );
  OAI2BB2XL U952 ( .B0(n1624), .B1(n1670), .A0N(\gbuff[19][4] ), .A1N(n1669), 
        .Y(n2183) );
  OAI2BB2XL U953 ( .B0(n1622), .B1(n1670), .A0N(\gbuff[19][5] ), .A1N(n1671), 
        .Y(n2182) );
  OAI2BB2XL U954 ( .B0(n1620), .B1(n1670), .A0N(\gbuff[19][6] ), .A1N(n1671), 
        .Y(n2181) );
  OAI2BB2XL U955 ( .B0(n1618), .B1(n1670), .A0N(\gbuff[19][7] ), .A1N(n1671), 
        .Y(n2180) );
  OAI2BB2XL U956 ( .B0(n1616), .B1(n1670), .A0N(\gbuff[19][8] ), .A1N(n1671), 
        .Y(n2179) );
  OAI2BB2XL U957 ( .B0(n1614), .B1(n1670), .A0N(\gbuff[19][9] ), .A1N(n1671), 
        .Y(n2178) );
  OAI2BB2XL U958 ( .B0(n1612), .B1(n1670), .A0N(\gbuff[19][10] ), .A1N(n1671), 
        .Y(n2177) );
  OAI2BB2XL U959 ( .B0(n1610), .B1(n1670), .A0N(\gbuff[19][11] ), .A1N(n1671), 
        .Y(n2176) );
  OAI2BB2XL U960 ( .B0(n1608), .B1(n1670), .A0N(\gbuff[19][12] ), .A1N(n1671), 
        .Y(n2175) );
  OAI2BB2XL U961 ( .B0(n1606), .B1(n1670), .A0N(\gbuff[19][13] ), .A1N(n1671), 
        .Y(n2174) );
  OAI2BB2XL U962 ( .B0(n1604), .B1(n1670), .A0N(\gbuff[19][14] ), .A1N(n1671), 
        .Y(n2173) );
  OAI2BB2XL U963 ( .B0(n1602), .B1(n1670), .A0N(\gbuff[19][15] ), .A1N(n1669), 
        .Y(n2172) );
  OAI2BB2XL U964 ( .B0(n1600), .B1(n1669), .A0N(\gbuff[19][16] ), .A1N(n1671), 
        .Y(n2171) );
  OAI2BB2XL U965 ( .B0(n1598), .B1(n1669), .A0N(\gbuff[19][17] ), .A1N(n1671), 
        .Y(n2170) );
  OAI2BB2XL U966 ( .B0(n1596), .B1(n2809), .A0N(\gbuff[19][18] ), .A1N(n1669), 
        .Y(n2169) );
  OAI2BB2XL U967 ( .B0(n1594), .B1(n1670), .A0N(\gbuff[19][19] ), .A1N(n1669), 
        .Y(n2168) );
  OAI2BB2XL U968 ( .B0(n1592), .B1(n2809), .A0N(\gbuff[19][20] ), .A1N(n1669), 
        .Y(n2167) );
  OAI2BB2XL U969 ( .B0(n1590), .B1(n2809), .A0N(\gbuff[19][21] ), .A1N(n1669), 
        .Y(n2166) );
  OAI2BB2XL U970 ( .B0(n1588), .B1(n1669), .A0N(\gbuff[19][22] ), .A1N(n1671), 
        .Y(n2165) );
  OAI2BB2XL U971 ( .B0(n1584), .B1(n2809), .A0N(\gbuff[19][24] ), .A1N(n1671), 
        .Y(n2163) );
  OAI2BB2XL U972 ( .B0(n1631), .B1(n1666), .A0N(\gbuff[20][0] ), .A1N(n1666), 
        .Y(n2155) );
  OAI2BB2XL U973 ( .B0(n1629), .B1(n1667), .A0N(\gbuff[20][1] ), .A1N(n1666), 
        .Y(n2154) );
  OAI2BB2XL U974 ( .B0(n1627), .B1(n1667), .A0N(\gbuff[20][2] ), .A1N(n1666), 
        .Y(n2153) );
  OAI2BB2XL U975 ( .B0(n1625), .B1(n1667), .A0N(\gbuff[20][3] ), .A1N(n1668), 
        .Y(n2152) );
  OAI2BB2XL U976 ( .B0(n1623), .B1(n1667), .A0N(\gbuff[20][4] ), .A1N(n1666), 
        .Y(n2151) );
  OAI2BB2XL U977 ( .B0(n1621), .B1(n1667), .A0N(\gbuff[20][5] ), .A1N(n1668), 
        .Y(n2150) );
  OAI2BB2XL U978 ( .B0(n1619), .B1(n1667), .A0N(\gbuff[20][6] ), .A1N(n1668), 
        .Y(n2149) );
  OAI2BB2XL U979 ( .B0(n1617), .B1(n1667), .A0N(\gbuff[20][7] ), .A1N(n1668), 
        .Y(n2148) );
  OAI2BB2XL U980 ( .B0(n1615), .B1(n1667), .A0N(\gbuff[20][8] ), .A1N(n1668), 
        .Y(n2147) );
  OAI2BB2XL U981 ( .B0(n1613), .B1(n1667), .A0N(\gbuff[20][9] ), .A1N(n1668), 
        .Y(n2146) );
  OAI2BB2XL U982 ( .B0(n1611), .B1(n1667), .A0N(\gbuff[20][10] ), .A1N(n1668), 
        .Y(n2145) );
  OAI2BB2XL U983 ( .B0(n1609), .B1(n1667), .A0N(\gbuff[20][11] ), .A1N(n1668), 
        .Y(n2144) );
  OAI2BB2XL U984 ( .B0(n1607), .B1(n1667), .A0N(\gbuff[20][12] ), .A1N(n1668), 
        .Y(n2143) );
  OAI2BB2XL U985 ( .B0(n1605), .B1(n2808), .A0N(\gbuff[20][13] ), .A1N(n1668), 
        .Y(n2142) );
  OAI2BB2XL U986 ( .B0(n1603), .B1(n2808), .A0N(\gbuff[20][14] ), .A1N(n1668), 
        .Y(n2141) );
  OAI2BB2XL U987 ( .B0(n1601), .B1(n2808), .A0N(\gbuff[20][15] ), .A1N(n1666), 
        .Y(n2140) );
  OAI2BB2XL U988 ( .B0(n1599), .B1(n1667), .A0N(\gbuff[20][16] ), .A1N(n1668), 
        .Y(n2139) );
  OAI2BB2XL U989 ( .B0(n1597), .B1(n1667), .A0N(\gbuff[20][17] ), .A1N(n1666), 
        .Y(n2138) );
  OAI2BB2XL U990 ( .B0(n1595), .B1(n1667), .A0N(\gbuff[20][18] ), .A1N(n1666), 
        .Y(n2137) );
  OAI2BB2XL U991 ( .B0(n1593), .B1(n2808), .A0N(\gbuff[20][19] ), .A1N(n1666), 
        .Y(n2136) );
  OAI2BB2XL U992 ( .B0(n1591), .B1(n1667), .A0N(\gbuff[20][20] ), .A1N(n1668), 
        .Y(n2135) );
  OAI2BB2XL U993 ( .B0(n1589), .B1(n1666), .A0N(\gbuff[20][21] ), .A1N(n1668), 
        .Y(n2134) );
  OAI2BB2XL U994 ( .B0(n1587), .B1(n2808), .A0N(\gbuff[20][22] ), .A1N(n1668), 
        .Y(n2133) );
  OAI2BB2XL U995 ( .B0(n1583), .B1(n1666), .A0N(\gbuff[20][24] ), .A1N(n1668), 
        .Y(n2131) );
  OAI2BB2XL U996 ( .B0(n1631), .B1(n1664), .A0N(\gbuff[21][0] ), .A1N(n1663), 
        .Y(n2123) );
  OAI2BB2XL U997 ( .B0(n1629), .B1(n1663), .A0N(\gbuff[21][1] ), .A1N(n1664), 
        .Y(n2122) );
  OAI2BB2XL U998 ( .B0(n1627), .B1(n1663), .A0N(\gbuff[21][2] ), .A1N(n1663), 
        .Y(n2121) );
  OAI2BB2XL U999 ( .B0(n1625), .B1(n1663), .A0N(\gbuff[21][3] ), .A1N(n1665), 
        .Y(n2120) );
  OAI2BB2XL U1000 ( .B0(n1623), .B1(n1663), .A0N(\gbuff[21][4] ), .A1N(n1664), 
        .Y(n2119) );
  OAI2BB2XL U1001 ( .B0(n1621), .B1(n1663), .A0N(\gbuff[21][5] ), .A1N(n1665), 
        .Y(n2118) );
  OAI2BB2XL U1002 ( .B0(n1619), .B1(n1663), .A0N(\gbuff[21][6] ), .A1N(n1665), 
        .Y(n2117) );
  OAI2BB2XL U1003 ( .B0(n1617), .B1(n1663), .A0N(\gbuff[21][7] ), .A1N(n1665), 
        .Y(n2116) );
  OAI2BB2XL U1004 ( .B0(n1615), .B1(n1663), .A0N(\gbuff[21][8] ), .A1N(n1665), 
        .Y(n2115) );
  OAI2BB2XL U1005 ( .B0(n1613), .B1(n1663), .A0N(\gbuff[21][9] ), .A1N(n1665), 
        .Y(n2114) );
  OAI2BB2XL U1006 ( .B0(n1611), .B1(n1663), .A0N(\gbuff[21][10] ), .A1N(n1665), 
        .Y(n2113) );
  OAI2BB2XL U1007 ( .B0(n1609), .B1(n1663), .A0N(\gbuff[21][11] ), .A1N(n1665), 
        .Y(n2112) );
  OAI2BB2XL U1008 ( .B0(n1607), .B1(n1663), .A0N(\gbuff[21][12] ), .A1N(n1665), 
        .Y(n2111) );
  OAI2BB2XL U1009 ( .B0(n1605), .B1(n1664), .A0N(\gbuff[21][13] ), .A1N(n1665), 
        .Y(n2110) );
  OAI2BB2XL U1010 ( .B0(n1603), .B1(n1664), .A0N(\gbuff[21][14] ), .A1N(n1665), 
        .Y(n2109) );
  OAI2BB2XL U1011 ( .B0(n1601), .B1(n1664), .A0N(\gbuff[21][15] ), .A1N(n1665), 
        .Y(n2108) );
  OAI2BB2XL U1012 ( .B0(n1599), .B1(n1664), .A0N(\gbuff[21][16] ), .A1N(n1665), 
        .Y(n2107) );
  OAI2BB2XL U1013 ( .B0(n1597), .B1(n1664), .A0N(\gbuff[21][17] ), .A1N(n1665), 
        .Y(n2106) );
  OAI2BB2XL U1014 ( .B0(n1595), .B1(n1664), .A0N(\gbuff[21][18] ), .A1N(n1663), 
        .Y(n2105) );
  OAI2BB2XL U1015 ( .B0(n1593), .B1(n1664), .A0N(\gbuff[21][19] ), .A1N(n1664), 
        .Y(n2104) );
  OAI2BB2XL U1016 ( .B0(n1591), .B1(n1664), .A0N(\gbuff[21][20] ), .A1N(n1665), 
        .Y(n2103) );
  OAI2BB2XL U1017 ( .B0(n1589), .B1(n1664), .A0N(\gbuff[21][21] ), .A1N(n1663), 
        .Y(n2102) );
  OAI2BB2XL U1018 ( .B0(n1587), .B1(n1664), .A0N(\gbuff[21][22] ), .A1N(n1665), 
        .Y(n2101) );
  OAI2BB2XL U1019 ( .B0(n1583), .B1(n1664), .A0N(\gbuff[21][24] ), .A1N(n1665), 
        .Y(n2099) );
  OAI2BB2XL U1020 ( .B0(n1631), .B1(n1661), .A0N(\gbuff[22][0] ), .A1N(n1660), 
        .Y(n2091) );
  OAI2BB2XL U1021 ( .B0(n1629), .B1(n1660), .A0N(\gbuff[22][1] ), .A1N(n1661), 
        .Y(n2090) );
  OAI2BB2XL U1022 ( .B0(n1627), .B1(n1660), .A0N(\gbuff[22][2] ), .A1N(n1660), 
        .Y(n2089) );
  OAI2BB2XL U1023 ( .B0(n1625), .B1(n1660), .A0N(\gbuff[22][3] ), .A1N(n1662), 
        .Y(n2088) );
  OAI2BB2XL U1024 ( .B0(n1623), .B1(n1660), .A0N(\gbuff[22][4] ), .A1N(n1661), 
        .Y(n2087) );
  OAI2BB2XL U1025 ( .B0(n1621), .B1(n1660), .A0N(\gbuff[22][5] ), .A1N(n1662), 
        .Y(n2086) );
  OAI2BB2XL U1026 ( .B0(n1619), .B1(n1660), .A0N(\gbuff[22][6] ), .A1N(n1662), 
        .Y(n2085) );
  OAI2BB2XL U1027 ( .B0(n1617), .B1(n1660), .A0N(\gbuff[22][7] ), .A1N(n1662), 
        .Y(n2084) );
  OAI2BB2XL U1028 ( .B0(n1615), .B1(n1660), .A0N(\gbuff[22][8] ), .A1N(n1662), 
        .Y(n2083) );
  OAI2BB2XL U1029 ( .B0(n1613), .B1(n1660), .A0N(\gbuff[22][9] ), .A1N(n1662), 
        .Y(n2082) );
  OAI2BB2XL U1030 ( .B0(n1611), .B1(n1660), .A0N(\gbuff[22][10] ), .A1N(n1662), 
        .Y(n2081) );
  OAI2BB2XL U1031 ( .B0(n1609), .B1(n1660), .A0N(\gbuff[22][11] ), .A1N(n1662), 
        .Y(n2080) );
  OAI2BB2XL U1032 ( .B0(n1607), .B1(n1660), .A0N(\gbuff[22][12] ), .A1N(n1662), 
        .Y(n2079) );
  OAI2BB2XL U1033 ( .B0(n1605), .B1(n1661), .A0N(\gbuff[22][13] ), .A1N(n1662), 
        .Y(n2078) );
  OAI2BB2XL U1034 ( .B0(n1603), .B1(n1661), .A0N(\gbuff[22][14] ), .A1N(n1662), 
        .Y(n2077) );
  OAI2BB2XL U1035 ( .B0(n1601), .B1(n1661), .A0N(\gbuff[22][15] ), .A1N(n1662), 
        .Y(n2076) );
  OAI2BB2XL U1036 ( .B0(n1599), .B1(n1661), .A0N(\gbuff[22][16] ), .A1N(n1662), 
        .Y(n2075) );
  OAI2BB2XL U1037 ( .B0(n1597), .B1(n1661), .A0N(\gbuff[22][17] ), .A1N(n1662), 
        .Y(n2074) );
  OAI2BB2XL U1038 ( .B0(n1595), .B1(n1661), .A0N(\gbuff[22][18] ), .A1N(n1660), 
        .Y(n2073) );
  OAI2BB2XL U1039 ( .B0(n1593), .B1(n1661), .A0N(\gbuff[22][19] ), .A1N(n1661), 
        .Y(n2072) );
  OAI2BB2XL U1040 ( .B0(n1591), .B1(n1661), .A0N(\gbuff[22][20] ), .A1N(n1662), 
        .Y(n2071) );
  OAI2BB2XL U1041 ( .B0(n1589), .B1(n1661), .A0N(\gbuff[22][21] ), .A1N(n1660), 
        .Y(n2070) );
  OAI2BB2XL U1042 ( .B0(n1587), .B1(n1661), .A0N(\gbuff[22][22] ), .A1N(n1662), 
        .Y(n2069) );
  OAI2BB2XL U1043 ( .B0(n1583), .B1(n1661), .A0N(\gbuff[22][24] ), .A1N(n1662), 
        .Y(n2067) );
  OAI2BB2XL U1044 ( .B0(n1631), .B1(n1658), .A0N(\gbuff[23][0] ), .A1N(n1657), 
        .Y(n2059) );
  OAI2BB2XL U1045 ( .B0(n1629), .B1(n1657), .A0N(\gbuff[23][1] ), .A1N(n1658), 
        .Y(n2058) );
  OAI2BB2XL U1046 ( .B0(n1627), .B1(n1657), .A0N(\gbuff[23][2] ), .A1N(n1657), 
        .Y(n2057) );
  OAI2BB2XL U1047 ( .B0(n1625), .B1(n1657), .A0N(\gbuff[23][3] ), .A1N(n1659), 
        .Y(n2056) );
  OAI2BB2XL U1048 ( .B0(n1623), .B1(n1657), .A0N(\gbuff[23][4] ), .A1N(n1658), 
        .Y(n2055) );
  OAI2BB2XL U1049 ( .B0(n1621), .B1(n1657), .A0N(\gbuff[23][5] ), .A1N(n1659), 
        .Y(n2054) );
  OAI2BB2XL U1050 ( .B0(n1619), .B1(n1657), .A0N(\gbuff[23][6] ), .A1N(n1659), 
        .Y(n2053) );
  OAI2BB2XL U1051 ( .B0(n1617), .B1(n1657), .A0N(\gbuff[23][7] ), .A1N(n1659), 
        .Y(n2052) );
  OAI2BB2XL U1052 ( .B0(n1615), .B1(n1657), .A0N(\gbuff[23][8] ), .A1N(n1659), 
        .Y(n2051) );
  OAI2BB2XL U1053 ( .B0(n1613), .B1(n1657), .A0N(\gbuff[23][9] ), .A1N(n1659), 
        .Y(n2050) );
  OAI2BB2XL U1054 ( .B0(n1611), .B1(n1657), .A0N(\gbuff[23][10] ), .A1N(n1659), 
        .Y(n2049) );
  OAI2BB2XL U1055 ( .B0(n1609), .B1(n1657), .A0N(\gbuff[23][11] ), .A1N(n1659), 
        .Y(n2048) );
  OAI2BB2XL U1056 ( .B0(n1607), .B1(n1657), .A0N(\gbuff[23][12] ), .A1N(n1659), 
        .Y(n2047) );
  OAI2BB2XL U1057 ( .B0(n1605), .B1(n1658), .A0N(\gbuff[23][13] ), .A1N(n1659), 
        .Y(n2046) );
  OAI2BB2XL U1058 ( .B0(n1603), .B1(n1658), .A0N(\gbuff[23][14] ), .A1N(n1659), 
        .Y(n2045) );
  OAI2BB2XL U1059 ( .B0(n1601), .B1(n1658), .A0N(\gbuff[23][15] ), .A1N(n1659), 
        .Y(n2044) );
  OAI2BB2XL U1060 ( .B0(n1599), .B1(n1658), .A0N(\gbuff[23][16] ), .A1N(n1659), 
        .Y(n2043) );
  OAI2BB2XL U1061 ( .B0(n1597), .B1(n1658), .A0N(\gbuff[23][17] ), .A1N(n1659), 
        .Y(n2042) );
  OAI2BB2XL U1062 ( .B0(n1595), .B1(n1658), .A0N(\gbuff[23][18] ), .A1N(n1657), 
        .Y(n2041) );
  OAI2BB2XL U1063 ( .B0(n1593), .B1(n1658), .A0N(\gbuff[23][19] ), .A1N(n1658), 
        .Y(n2040) );
  OAI2BB2XL U1064 ( .B0(n1591), .B1(n1658), .A0N(\gbuff[23][20] ), .A1N(n1659), 
        .Y(n2039) );
  OAI2BB2XL U1065 ( .B0(n1589), .B1(n1658), .A0N(\gbuff[23][21] ), .A1N(n1657), 
        .Y(n2038) );
  OAI2BB2XL U1066 ( .B0(n1587), .B1(n1658), .A0N(\gbuff[23][22] ), .A1N(n1659), 
        .Y(n2037) );
  OAI2BB2XL U1067 ( .B0(n1583), .B1(n1658), .A0N(\gbuff[23][24] ), .A1N(n1659), 
        .Y(n2035) );
  OAI2BB2XL U1068 ( .B0(n1631), .B1(n1655), .A0N(\gbuff[24][0] ), .A1N(n1654), 
        .Y(n2027) );
  OAI2BB2XL U1069 ( .B0(n1629), .B1(n1655), .A0N(\gbuff[24][1] ), .A1N(n1654), 
        .Y(n2026) );
  OAI2BB2XL U1070 ( .B0(n1627), .B1(n1655), .A0N(\gbuff[24][2] ), .A1N(n1654), 
        .Y(n2025) );
  OAI2BB2XL U1071 ( .B0(n1625), .B1(n1655), .A0N(\gbuff[24][3] ), .A1N(n1656), 
        .Y(n2024) );
  OAI2BB2XL U1072 ( .B0(n1623), .B1(n1655), .A0N(\gbuff[24][4] ), .A1N(n1654), 
        .Y(n2023) );
  OAI2BB2XL U1073 ( .B0(n1621), .B1(n1655), .A0N(\gbuff[24][5] ), .A1N(n1656), 
        .Y(n2022) );
  OAI2BB2XL U1074 ( .B0(n1619), .B1(n1655), .A0N(\gbuff[24][6] ), .A1N(n1656), 
        .Y(n2021) );
  OAI2BB2XL U1075 ( .B0(n1617), .B1(n1655), .A0N(\gbuff[24][7] ), .A1N(n1656), 
        .Y(n2020) );
  OAI2BB2XL U1076 ( .B0(n1615), .B1(n1655), .A0N(\gbuff[24][8] ), .A1N(n1656), 
        .Y(n2019) );
  OAI2BB2XL U1077 ( .B0(n1613), .B1(n1655), .A0N(\gbuff[24][9] ), .A1N(n1656), 
        .Y(n2018) );
  OAI2BB2XL U1078 ( .B0(n1611), .B1(n1655), .A0N(\gbuff[24][10] ), .A1N(n1656), 
        .Y(n2017) );
  OAI2BB2XL U1079 ( .B0(n1609), .B1(n1655), .A0N(\gbuff[24][11] ), .A1N(n1656), 
        .Y(n2016) );
  OAI2BB2XL U1080 ( .B0(n1607), .B1(n1655), .A0N(\gbuff[24][12] ), .A1N(n1656), 
        .Y(n2015) );
  OAI2BB2XL U1081 ( .B0(n1605), .B1(n1655), .A0N(\gbuff[24][13] ), .A1N(n1656), 
        .Y(n2014) );
  OAI2BB2XL U1082 ( .B0(n1603), .B1(n1655), .A0N(\gbuff[24][14] ), .A1N(n1656), 
        .Y(n2013) );
  OAI2BB2XL U1083 ( .B0(n1601), .B1(n1655), .A0N(\gbuff[24][15] ), .A1N(n1654), 
        .Y(n2012) );
  OAI2BB2XL U1084 ( .B0(n1599), .B1(n1654), .A0N(\gbuff[24][16] ), .A1N(n1656), 
        .Y(n2011) );
  OAI2BB2XL U1085 ( .B0(n1597), .B1(n1654), .A0N(\gbuff[24][17] ), .A1N(n1656), 
        .Y(n2010) );
  OAI2BB2XL U1086 ( .B0(n1595), .B1(n2804), .A0N(\gbuff[24][18] ), .A1N(n1654), 
        .Y(n2009) );
  OAI2BB2XL U1087 ( .B0(n1593), .B1(n1655), .A0N(\gbuff[24][19] ), .A1N(n1654), 
        .Y(n2008) );
  OAI2BB2XL U1088 ( .B0(n1591), .B1(n2804), .A0N(\gbuff[24][20] ), .A1N(n1654), 
        .Y(n2007) );
  OAI2BB2XL U1089 ( .B0(n1589), .B1(n2804), .A0N(\gbuff[24][21] ), .A1N(n1654), 
        .Y(n2006) );
  OAI2BB2XL U1090 ( .B0(n1587), .B1(n1654), .A0N(\gbuff[24][22] ), .A1N(n1656), 
        .Y(n2005) );
  OAI2BB2XL U1091 ( .B0(n1583), .B1(n2804), .A0N(\gbuff[24][24] ), .A1N(n1656), 
        .Y(n2003) );
  OAI2BB2XL U1092 ( .B0(n1631), .B1(n1652), .A0N(\gbuff[25][0] ), .A1N(n1651), 
        .Y(n1995) );
  OAI2BB2XL U1093 ( .B0(n1629), .B1(n1652), .A0N(\gbuff[25][1] ), .A1N(n1651), 
        .Y(n1994) );
  OAI2BB2XL U1094 ( .B0(n1627), .B1(n1652), .A0N(\gbuff[25][2] ), .A1N(n1651), 
        .Y(n1993) );
  OAI2BB2XL U1095 ( .B0(n1625), .B1(n1652), .A0N(\gbuff[25][3] ), .A1N(n1653), 
        .Y(n1992) );
  OAI2BB2XL U1096 ( .B0(n1623), .B1(n1652), .A0N(\gbuff[25][4] ), .A1N(n1651), 
        .Y(n1991) );
  OAI2BB2XL U1097 ( .B0(n1621), .B1(n1652), .A0N(\gbuff[25][5] ), .A1N(n1653), 
        .Y(n1990) );
  OAI2BB2XL U1098 ( .B0(n1619), .B1(n1652), .A0N(\gbuff[25][6] ), .A1N(n1653), 
        .Y(n1989) );
  OAI2BB2XL U1099 ( .B0(n1617), .B1(n1652), .A0N(\gbuff[25][7] ), .A1N(n1653), 
        .Y(n1988) );
  OAI2BB2XL U1100 ( .B0(n1615), .B1(n1652), .A0N(\gbuff[25][8] ), .A1N(n1653), 
        .Y(n1987) );
  OAI2BB2XL U1101 ( .B0(n1613), .B1(n1652), .A0N(\gbuff[25][9] ), .A1N(n1653), 
        .Y(n1986) );
  OAI2BB2XL U1102 ( .B0(n1611), .B1(n1652), .A0N(\gbuff[25][10] ), .A1N(n1653), 
        .Y(n1985) );
  OAI2BB2XL U1103 ( .B0(n1609), .B1(n1652), .A0N(\gbuff[25][11] ), .A1N(n1653), 
        .Y(n1984) );
  OAI2BB2XL U1104 ( .B0(n1607), .B1(n1652), .A0N(\gbuff[25][12] ), .A1N(n1653), 
        .Y(n1983) );
  OAI2BB2XL U1105 ( .B0(n1605), .B1(n1652), .A0N(\gbuff[25][13] ), .A1N(n1653), 
        .Y(n1982) );
  OAI2BB2XL U1106 ( .B0(n1603), .B1(n1652), .A0N(\gbuff[25][14] ), .A1N(n1653), 
        .Y(n1981) );
  OAI2BB2XL U1107 ( .B0(n1601), .B1(n1652), .A0N(\gbuff[25][15] ), .A1N(n1651), 
        .Y(n1980) );
  OAI2BB2XL U1108 ( .B0(n1599), .B1(n1651), .A0N(\gbuff[25][16] ), .A1N(n1653), 
        .Y(n1979) );
  OAI2BB2XL U1109 ( .B0(n1597), .B1(n1651), .A0N(\gbuff[25][17] ), .A1N(n1653), 
        .Y(n1978) );
  OAI2BB2XL U1110 ( .B0(n1595), .B1(n2802), .A0N(\gbuff[25][18] ), .A1N(n1651), 
        .Y(n1977) );
  OAI2BB2XL U1111 ( .B0(n1593), .B1(n1652), .A0N(\gbuff[25][19] ), .A1N(n1651), 
        .Y(n1976) );
  OAI2BB2XL U1112 ( .B0(n1591), .B1(n2802), .A0N(\gbuff[25][20] ), .A1N(n1651), 
        .Y(n1975) );
  OAI2BB2XL U1113 ( .B0(n1589), .B1(n2802), .A0N(\gbuff[25][21] ), .A1N(n1651), 
        .Y(n1974) );
  OAI2BB2XL U1114 ( .B0(n1587), .B1(n1651), .A0N(\gbuff[25][22] ), .A1N(n1653), 
        .Y(n1973) );
  OAI2BB2XL U1115 ( .B0(n1583), .B1(n2802), .A0N(\gbuff[25][24] ), .A1N(n1653), 
        .Y(n1971) );
  OAI2BB2XL U1116 ( .B0(n1631), .B1(n1649), .A0N(\gbuff[26][0] ), .A1N(n1648), 
        .Y(n1963) );
  OAI2BB2XL U1117 ( .B0(n1629), .B1(n1649), .A0N(\gbuff[26][1] ), .A1N(n1648), 
        .Y(n1962) );
  OAI2BB2XL U1118 ( .B0(n1627), .B1(n1649), .A0N(\gbuff[26][2] ), .A1N(n1648), 
        .Y(n1961) );
  OAI2BB2XL U1119 ( .B0(n1625), .B1(n1649), .A0N(\gbuff[26][3] ), .A1N(n1650), 
        .Y(n1960) );
  OAI2BB2XL U1120 ( .B0(n1623), .B1(n1649), .A0N(\gbuff[26][4] ), .A1N(n1648), 
        .Y(n1959) );
  OAI2BB2XL U1121 ( .B0(n1621), .B1(n1649), .A0N(\gbuff[26][5] ), .A1N(n1650), 
        .Y(n1958) );
  OAI2BB2XL U1122 ( .B0(n1619), .B1(n1649), .A0N(\gbuff[26][6] ), .A1N(n1650), 
        .Y(n1957) );
  OAI2BB2XL U1123 ( .B0(n1617), .B1(n1649), .A0N(\gbuff[26][7] ), .A1N(n1650), 
        .Y(n1956) );
  OAI2BB2XL U1124 ( .B0(n1615), .B1(n1649), .A0N(\gbuff[26][8] ), .A1N(n1650), 
        .Y(n1955) );
  OAI2BB2XL U1125 ( .B0(n1613), .B1(n1649), .A0N(\gbuff[26][9] ), .A1N(n1650), 
        .Y(n1954) );
  OAI2BB2XL U1126 ( .B0(n1611), .B1(n1649), .A0N(\gbuff[26][10] ), .A1N(n1650), 
        .Y(n1953) );
  OAI2BB2XL U1127 ( .B0(n1609), .B1(n1649), .A0N(\gbuff[26][11] ), .A1N(n1650), 
        .Y(n1952) );
  OAI2BB2XL U1128 ( .B0(n1607), .B1(n1649), .A0N(\gbuff[26][12] ), .A1N(n1650), 
        .Y(n1951) );
  OAI2BB2XL U1129 ( .B0(n1605), .B1(n1649), .A0N(\gbuff[26][13] ), .A1N(n1650), 
        .Y(n1950) );
  OAI2BB2XL U1130 ( .B0(n1603), .B1(n1649), .A0N(\gbuff[26][14] ), .A1N(n1650), 
        .Y(n1949) );
  OAI2BB2XL U1131 ( .B0(n1601), .B1(n1649), .A0N(\gbuff[26][15] ), .A1N(n1648), 
        .Y(n1948) );
  OAI2BB2XL U1132 ( .B0(n1599), .B1(n1648), .A0N(\gbuff[26][16] ), .A1N(n1650), 
        .Y(n1947) );
  OAI2BB2XL U1133 ( .B0(n1597), .B1(n1648), .A0N(\gbuff[26][17] ), .A1N(n1650), 
        .Y(n1946) );
  OAI2BB2XL U1134 ( .B0(n1595), .B1(n2801), .A0N(\gbuff[26][18] ), .A1N(n1648), 
        .Y(n1945) );
  OAI2BB2XL U1135 ( .B0(n1593), .B1(n1649), .A0N(\gbuff[26][19] ), .A1N(n1648), 
        .Y(n1944) );
  OAI2BB2XL U1136 ( .B0(n1591), .B1(n2801), .A0N(\gbuff[26][20] ), .A1N(n1648), 
        .Y(n1943) );
  OAI2BB2XL U1137 ( .B0(n1589), .B1(n2801), .A0N(\gbuff[26][21] ), .A1N(n1648), 
        .Y(n1942) );
  OAI2BB2XL U1138 ( .B0(n1587), .B1(n1648), .A0N(\gbuff[26][22] ), .A1N(n1650), 
        .Y(n1941) );
  OAI2BB2XL U1139 ( .B0(n1583), .B1(n2801), .A0N(\gbuff[26][24] ), .A1N(n1650), 
        .Y(n1939) );
  OAI2BB2XL U1140 ( .B0(n1631), .B1(n1646), .A0N(\gbuff[27][0] ), .A1N(n1645), 
        .Y(n1931) );
  OAI2BB2XL U1141 ( .B0(n1629), .B1(n1646), .A0N(\gbuff[27][1] ), .A1N(n1645), 
        .Y(n1930) );
  OAI2BB2XL U1142 ( .B0(n1627), .B1(n1646), .A0N(\gbuff[27][2] ), .A1N(n1645), 
        .Y(n1929) );
  OAI2BB2XL U1143 ( .B0(n1625), .B1(n1646), .A0N(\gbuff[27][3] ), .A1N(n1647), 
        .Y(n1928) );
  OAI2BB2XL U1144 ( .B0(n1623), .B1(n1646), .A0N(\gbuff[27][4] ), .A1N(n1645), 
        .Y(n1927) );
  OAI2BB2XL U1145 ( .B0(n1621), .B1(n1646), .A0N(\gbuff[27][5] ), .A1N(n1647), 
        .Y(n1926) );
  OAI2BB2XL U1146 ( .B0(n1619), .B1(n1646), .A0N(\gbuff[27][6] ), .A1N(n1647), 
        .Y(n1925) );
  OAI2BB2XL U1147 ( .B0(n1617), .B1(n1646), .A0N(\gbuff[27][7] ), .A1N(n1647), 
        .Y(n1924) );
  OAI2BB2XL U1148 ( .B0(n1615), .B1(n1646), .A0N(\gbuff[27][8] ), .A1N(n1647), 
        .Y(n1923) );
  OAI2BB2XL U1149 ( .B0(n1613), .B1(n1646), .A0N(\gbuff[27][9] ), .A1N(n1647), 
        .Y(n1922) );
  OAI2BB2XL U1150 ( .B0(n1611), .B1(n1646), .A0N(\gbuff[27][10] ), .A1N(n1647), 
        .Y(n1921) );
  OAI2BB2XL U1151 ( .B0(n1609), .B1(n1646), .A0N(\gbuff[27][11] ), .A1N(n1647), 
        .Y(n1920) );
  OAI2BB2XL U1152 ( .B0(n1607), .B1(n1646), .A0N(\gbuff[27][12] ), .A1N(n1647), 
        .Y(n1919) );
  OAI2BB2XL U1153 ( .B0(n1605), .B1(n1646), .A0N(\gbuff[27][13] ), .A1N(n1647), 
        .Y(n1918) );
  OAI2BB2XL U1154 ( .B0(n1603), .B1(n1646), .A0N(\gbuff[27][14] ), .A1N(n1647), 
        .Y(n1917) );
  OAI2BB2XL U1155 ( .B0(n1601), .B1(n1646), .A0N(\gbuff[27][15] ), .A1N(n1645), 
        .Y(n1916) );
  OAI2BB2XL U1156 ( .B0(n1599), .B1(n1645), .A0N(\gbuff[27][16] ), .A1N(n1647), 
        .Y(n1915) );
  OAI2BB2XL U1157 ( .B0(n1597), .B1(n2800), .A0N(\gbuff[27][17] ), .A1N(n1645), 
        .Y(n1914) );
  OAI2BB2XL U1158 ( .B0(n1595), .B1(n2800), .A0N(\gbuff[27][18] ), .A1N(n1645), 
        .Y(n1913) );
  OAI2BB2XL U1159 ( .B0(n1593), .B1(n1646), .A0N(\gbuff[27][19] ), .A1N(n1645), 
        .Y(n1912) );
  OAI2BB2XL U1160 ( .B0(n1591), .B1(n2800), .A0N(\gbuff[27][20] ), .A1N(n1645), 
        .Y(n1911) );
  OAI2BB2XL U1161 ( .B0(n1589), .B1(n2800), .A0N(\gbuff[27][21] ), .A1N(n1645), 
        .Y(n1910) );
  OAI2BB2XL U1162 ( .B0(n1587), .B1(n1645), .A0N(\gbuff[27][22] ), .A1N(n1647), 
        .Y(n1909) );
  OAI2BB2XL U1163 ( .B0(n1583), .B1(n2800), .A0N(\gbuff[27][24] ), .A1N(n1647), 
        .Y(n1907) );
  OAI2BB2XL U1164 ( .B0(n1631), .B1(n1642), .A0N(\gbuff[28][0] ), .A1N(n1643), 
        .Y(n1899) );
  OAI2BB2XL U1165 ( .B0(n1629), .B1(n1642), .A0N(\gbuff[28][1] ), .A1N(n1644), 
        .Y(n1898) );
  OAI2BB2XL U1166 ( .B0(n1627), .B1(n1642), .A0N(\gbuff[28][2] ), .A1N(n1643), 
        .Y(n1897) );
  OAI2BB2XL U1167 ( .B0(n1625), .B1(n1642), .A0N(\gbuff[28][3] ), .A1N(n1644), 
        .Y(n1896) );
  OAI2BB2XL U1168 ( .B0(n1623), .B1(n1642), .A0N(\gbuff[28][4] ), .A1N(n1644), 
        .Y(n1895) );
  OAI2BB2XL U1169 ( .B0(n1621), .B1(n1642), .A0N(\gbuff[28][5] ), .A1N(n1644), 
        .Y(n1894) );
  OAI2BB2XL U1170 ( .B0(n1619), .B1(n1642), .A0N(\gbuff[28][6] ), .A1N(n1644), 
        .Y(n1893) );
  OAI2BB2XL U1171 ( .B0(n1617), .B1(n1642), .A0N(\gbuff[28][7] ), .A1N(n1644), 
        .Y(n1892) );
  OAI2BB2XL U1172 ( .B0(n1615), .B1(n1642), .A0N(\gbuff[28][8] ), .A1N(n1644), 
        .Y(n1891) );
  OAI2BB2XL U1173 ( .B0(n1613), .B1(n1642), .A0N(\gbuff[28][9] ), .A1N(n1644), 
        .Y(n1890) );
  OAI2BB2XL U1174 ( .B0(n1611), .B1(n1642), .A0N(\gbuff[28][10] ), .A1N(n1644), 
        .Y(n1889) );
  OAI2BB2XL U1175 ( .B0(n1609), .B1(n1642), .A0N(\gbuff[28][11] ), .A1N(n1644), 
        .Y(n1888) );
  OAI2BB2XL U1176 ( .B0(n1607), .B1(n1642), .A0N(\gbuff[28][12] ), .A1N(n1644), 
        .Y(n1887) );
  OAI2BB2XL U1177 ( .B0(n1605), .B1(n1642), .A0N(\gbuff[28][13] ), .A1N(n1644), 
        .Y(n1886) );
  OAI2BB2XL U1178 ( .B0(n1603), .B1(n1642), .A0N(\gbuff[28][14] ), .A1N(n1644), 
        .Y(n1885) );
  OAI2BB2XL U1179 ( .B0(n1601), .B1(n1642), .A0N(\gbuff[28][15] ), .A1N(n1643), 
        .Y(n1884) );
  OAI2BB2XL U1180 ( .B0(n1599), .B1(n1642), .A0N(\gbuff[28][16] ), .A1N(n1644), 
        .Y(n1883) );
  OAI2BB2XL U1181 ( .B0(n1597), .B1(n1642), .A0N(\gbuff[28][17] ), .A1N(n1643), 
        .Y(n1882) );
  OAI2BB2XL U1182 ( .B0(n1595), .B1(n1643), .A0N(\gbuff[28][18] ), .A1N(n1643), 
        .Y(n1881) );
  OAI2BB2XL U1183 ( .B0(n1593), .B1(n1642), .A0N(\gbuff[28][19] ), .A1N(n1643), 
        .Y(n1880) );
  OAI2BB2XL U1184 ( .B0(n1591), .B1(n1642), .A0N(\gbuff[28][20] ), .A1N(n1643), 
        .Y(n1879) );
  OAI2BB2XL U1185 ( .B0(n1589), .B1(n1643), .A0N(\gbuff[28][21] ), .A1N(n1643), 
        .Y(n1878) );
  OAI2BB2XL U1186 ( .B0(n1587), .B1(n1642), .A0N(\gbuff[28][22] ), .A1N(n1644), 
        .Y(n1877) );
  OAI2BB2XL U1187 ( .B0(n1583), .B1(n1643), .A0N(\gbuff[28][24] ), .A1N(n1644), 
        .Y(n1875) );
  OAI2BB2XL U1188 ( .B0(n1631), .B1(n1639), .A0N(\gbuff[29][0] ), .A1N(n1640), 
        .Y(n1867) );
  OAI2BB2XL U1189 ( .B0(n1629), .B1(n1639), .A0N(\gbuff[29][1] ), .A1N(n1641), 
        .Y(n1866) );
  OAI2BB2XL U1190 ( .B0(n1627), .B1(n1639), .A0N(\gbuff[29][2] ), .A1N(n1640), 
        .Y(n1865) );
  OAI2BB2XL U1191 ( .B0(n1625), .B1(n1639), .A0N(\gbuff[29][3] ), .A1N(n1641), 
        .Y(n1864) );
  OAI2BB2XL U1192 ( .B0(n1623), .B1(n1639), .A0N(\gbuff[29][4] ), .A1N(n1641), 
        .Y(n1863) );
  OAI2BB2XL U1193 ( .B0(n1621), .B1(n1639), .A0N(\gbuff[29][5] ), .A1N(n1641), 
        .Y(n1862) );
  OAI2BB2XL U1194 ( .B0(n1619), .B1(n1639), .A0N(\gbuff[29][6] ), .A1N(n1641), 
        .Y(n1861) );
  OAI2BB2XL U1195 ( .B0(n1617), .B1(n1639), .A0N(\gbuff[29][7] ), .A1N(n1641), 
        .Y(n1860) );
  OAI2BB2XL U1196 ( .B0(n1615), .B1(n1639), .A0N(\gbuff[29][8] ), .A1N(n1641), 
        .Y(n1859) );
  OAI2BB2XL U1197 ( .B0(n1613), .B1(n1639), .A0N(\gbuff[29][9] ), .A1N(n1641), 
        .Y(n1858) );
  OAI2BB2XL U1198 ( .B0(n1611), .B1(n1639), .A0N(\gbuff[29][10] ), .A1N(n1641), 
        .Y(n1857) );
  OAI2BB2XL U1199 ( .B0(n1609), .B1(n1639), .A0N(\gbuff[29][11] ), .A1N(n1641), 
        .Y(n1856) );
  OAI2BB2XL U1200 ( .B0(n1607), .B1(n1639), .A0N(\gbuff[29][12] ), .A1N(n1641), 
        .Y(n1855) );
  OAI2BB2XL U1201 ( .B0(n1605), .B1(n1639), .A0N(\gbuff[29][13] ), .A1N(n1641), 
        .Y(n1854) );
  OAI2BB2XL U1202 ( .B0(n1603), .B1(n1639), .A0N(\gbuff[29][14] ), .A1N(n1641), 
        .Y(n1853) );
  OAI2BB2XL U1203 ( .B0(n1601), .B1(n1639), .A0N(\gbuff[29][15] ), .A1N(n1640), 
        .Y(n1852) );
  OAI2BB2XL U1204 ( .B0(n1599), .B1(n1639), .A0N(\gbuff[29][16] ), .A1N(n1641), 
        .Y(n1851) );
  OAI2BB2XL U1205 ( .B0(n1597), .B1(n1639), .A0N(\gbuff[29][17] ), .A1N(n1640), 
        .Y(n1850) );
  OAI2BB2XL U1206 ( .B0(n1595), .B1(n1640), .A0N(\gbuff[29][18] ), .A1N(n1640), 
        .Y(n1849) );
  OAI2BB2XL U1207 ( .B0(n1593), .B1(n1639), .A0N(\gbuff[29][19] ), .A1N(n1640), 
        .Y(n1848) );
  OAI2BB2XL U1208 ( .B0(n1591), .B1(n1639), .A0N(\gbuff[29][20] ), .A1N(n1640), 
        .Y(n1847) );
  OAI2BB2XL U1209 ( .B0(n1589), .B1(n1640), .A0N(\gbuff[29][21] ), .A1N(n1640), 
        .Y(n1846) );
  OAI2BB2XL U1210 ( .B0(n1587), .B1(n1639), .A0N(\gbuff[29][22] ), .A1N(n1641), 
        .Y(n1845) );
  OAI2BB2XL U1211 ( .B0(n1583), .B1(n1640), .A0N(\gbuff[29][24] ), .A1N(n1641), 
        .Y(n1843) );
  OAI2BB2XL U1212 ( .B0(n1631), .B1(n1636), .A0N(\gbuff[30][0] ), .A1N(n1637), 
        .Y(n1835) );
  OAI2BB2XL U1213 ( .B0(n1629), .B1(n1636), .A0N(\gbuff[30][1] ), .A1N(n1638), 
        .Y(n1834) );
  OAI2BB2XL U1214 ( .B0(n1627), .B1(n1636), .A0N(\gbuff[30][2] ), .A1N(n1637), 
        .Y(n1833) );
  OAI2BB2XL U1215 ( .B0(n1625), .B1(n1636), .A0N(\gbuff[30][3] ), .A1N(n1638), 
        .Y(n1832) );
  OAI2BB2XL U1216 ( .B0(n1623), .B1(n1636), .A0N(\gbuff[30][4] ), .A1N(n1638), 
        .Y(n1831) );
  OAI2BB2XL U1217 ( .B0(n1621), .B1(n1636), .A0N(\gbuff[30][5] ), .A1N(n1638), 
        .Y(n1830) );
  OAI2BB2XL U1218 ( .B0(n1619), .B1(n1636), .A0N(\gbuff[30][6] ), .A1N(n1638), 
        .Y(n1829) );
  OAI2BB2XL U1219 ( .B0(n1617), .B1(n1636), .A0N(\gbuff[30][7] ), .A1N(n1638), 
        .Y(n1828) );
  OAI2BB2XL U1220 ( .B0(n1615), .B1(n1636), .A0N(\gbuff[30][8] ), .A1N(n1638), 
        .Y(n1827) );
  OAI2BB2XL U1221 ( .B0(n1613), .B1(n1636), .A0N(\gbuff[30][9] ), .A1N(n1638), 
        .Y(n1826) );
  OAI2BB2XL U1222 ( .B0(n1611), .B1(n1636), .A0N(\gbuff[30][10] ), .A1N(n1638), 
        .Y(n1825) );
  OAI2BB2XL U1223 ( .B0(n1609), .B1(n1636), .A0N(\gbuff[30][11] ), .A1N(n1638), 
        .Y(n1824) );
  OAI2BB2XL U1224 ( .B0(n1607), .B1(n1636), .A0N(\gbuff[30][12] ), .A1N(n1638), 
        .Y(n1823) );
  OAI2BB2XL U1225 ( .B0(n1605), .B1(n1636), .A0N(\gbuff[30][13] ), .A1N(n1638), 
        .Y(n1822) );
  OAI2BB2XL U1226 ( .B0(n1603), .B1(n1636), .A0N(\gbuff[30][14] ), .A1N(n1638), 
        .Y(n1821) );
  OAI2BB2XL U1227 ( .B0(n1601), .B1(n1636), .A0N(\gbuff[30][15] ), .A1N(n1637), 
        .Y(n1820) );
  OAI2BB2XL U1228 ( .B0(n1599), .B1(n1636), .A0N(\gbuff[30][16] ), .A1N(n1638), 
        .Y(n1819) );
  OAI2BB2XL U1229 ( .B0(n1597), .B1(n1636), .A0N(\gbuff[30][17] ), .A1N(n1637), 
        .Y(n1818) );
  OAI2BB2XL U1230 ( .B0(n1595), .B1(n1637), .A0N(\gbuff[30][18] ), .A1N(n1637), 
        .Y(n1817) );
  OAI2BB2XL U1231 ( .B0(n1593), .B1(n1636), .A0N(\gbuff[30][19] ), .A1N(n1637), 
        .Y(n1816) );
  OAI2BB2XL U1232 ( .B0(n1591), .B1(n1636), .A0N(\gbuff[30][20] ), .A1N(n1637), 
        .Y(n1815) );
  OAI2BB2XL U1233 ( .B0(n1589), .B1(n1637), .A0N(\gbuff[30][21] ), .A1N(n1637), 
        .Y(n1814) );
  OAI2BB2XL U1234 ( .B0(n1587), .B1(n1636), .A0N(\gbuff[30][22] ), .A1N(n1638), 
        .Y(n1813) );
  OAI2BB2XL U1235 ( .B0(n1583), .B1(n1637), .A0N(\gbuff[30][24] ), .A1N(n1638), 
        .Y(n1811) );
  OAI2BB2XL U1236 ( .B0(n1631), .B1(n1633), .A0N(\gbuff[31][0] ), .A1N(n1634), 
        .Y(n1803) );
  OAI2BB2XL U1237 ( .B0(n1629), .B1(n1633), .A0N(\gbuff[31][1] ), .A1N(n1635), 
        .Y(n1802) );
  OAI2BB2XL U1238 ( .B0(n1627), .B1(n1633), .A0N(\gbuff[31][2] ), .A1N(n1634), 
        .Y(n1801) );
  OAI2BB2XL U1239 ( .B0(n1625), .B1(n1633), .A0N(\gbuff[31][3] ), .A1N(n1635), 
        .Y(n1800) );
  OAI2BB2XL U1240 ( .B0(n1623), .B1(n1633), .A0N(\gbuff[31][4] ), .A1N(n1635), 
        .Y(n1799) );
  OAI2BB2XL U1241 ( .B0(n1621), .B1(n1633), .A0N(\gbuff[31][5] ), .A1N(n1635), 
        .Y(n1798) );
  OAI2BB2XL U1242 ( .B0(n1619), .B1(n1633), .A0N(\gbuff[31][6] ), .A1N(n1635), 
        .Y(n1797) );
  OAI2BB2XL U1243 ( .B0(n1617), .B1(n1633), .A0N(\gbuff[31][7] ), .A1N(n1635), 
        .Y(n1796) );
  OAI2BB2XL U1244 ( .B0(n1615), .B1(n1633), .A0N(\gbuff[31][8] ), .A1N(n1635), 
        .Y(n1795) );
  OAI2BB2XL U1245 ( .B0(n1613), .B1(n1633), .A0N(\gbuff[31][9] ), .A1N(n1635), 
        .Y(n1794) );
  OAI2BB2XL U1246 ( .B0(n1611), .B1(n1633), .A0N(\gbuff[31][10] ), .A1N(n1635), 
        .Y(n1793) );
  OAI2BB2XL U1247 ( .B0(n1609), .B1(n1633), .A0N(\gbuff[31][11] ), .A1N(n1635), 
        .Y(n1792) );
  OAI2BB2XL U1248 ( .B0(n1607), .B1(n1633), .A0N(\gbuff[31][12] ), .A1N(n1635), 
        .Y(n1791) );
  OAI2BB2XL U1249 ( .B0(n1605), .B1(n1633), .A0N(\gbuff[31][13] ), .A1N(n1635), 
        .Y(n1790) );
  OAI2BB2XL U1250 ( .B0(n1603), .B1(n1633), .A0N(\gbuff[31][14] ), .A1N(n1635), 
        .Y(n1789) );
  OAI2BB2XL U1251 ( .B0(n1601), .B1(n1633), .A0N(\gbuff[31][15] ), .A1N(n1634), 
        .Y(n1788) );
  OAI2BB2XL U1252 ( .B0(n1599), .B1(n1633), .A0N(\gbuff[31][16] ), .A1N(n1635), 
        .Y(n1787) );
  OAI2BB2XL U1253 ( .B0(n1597), .B1(n1633), .A0N(\gbuff[31][17] ), .A1N(n1634), 
        .Y(n1786) );
  OAI2BB2XL U1254 ( .B0(n1595), .B1(n1634), .A0N(\gbuff[31][18] ), .A1N(n1634), 
        .Y(n1785) );
  OAI2BB2XL U1255 ( .B0(n1593), .B1(n1633), .A0N(\gbuff[31][19] ), .A1N(n1634), 
        .Y(n1784) );
  OAI2BB2XL U1256 ( .B0(n1591), .B1(n1633), .A0N(\gbuff[31][20] ), .A1N(n1634), 
        .Y(n1783) );
  OAI2BB2XL U1257 ( .B0(n1589), .B1(n1634), .A0N(\gbuff[31][21] ), .A1N(n1634), 
        .Y(n1782) );
  OAI2BB2XL U1258 ( .B0(n1587), .B1(n1633), .A0N(\gbuff[31][22] ), .A1N(n1635), 
        .Y(n1781) );
  OAI2BB2XL U1259 ( .B0(n1583), .B1(n1634), .A0N(\gbuff[31][24] ), .A1N(n1635), 
        .Y(n1779) );
  OAI2BB2XL U1260 ( .B0(n1726), .B1(n1771), .A0N(\gbuff[0][0] ), .A1N(n1), .Y(
        n2795) );
  OAI2BB2XL U1261 ( .B0(n1726), .B1(n1770), .A0N(\gbuff[0][1] ), .A1N(n1), .Y(
        n2794) );
  OAI2BB2XL U1262 ( .B0(n1726), .B1(n1769), .A0N(\gbuff[0][2] ), .A1N(n1), .Y(
        n2793) );
  OAI2BB2XL U1263 ( .B0(n1726), .B1(n1768), .A0N(\gbuff[0][3] ), .A1N(n1728), 
        .Y(n2792) );
  OAI2BB2XL U1264 ( .B0(n1726), .B1(n1767), .A0N(\gbuff[0][4] ), .A1N(n1728), 
        .Y(n2791) );
  OAI2BB2XL U1265 ( .B0(n1726), .B1(n1766), .A0N(\gbuff[0][5] ), .A1N(n1728), 
        .Y(n2790) );
  OAI2BB2XL U1266 ( .B0(n1726), .B1(n1765), .A0N(\gbuff[0][6] ), .A1N(n1728), 
        .Y(n2789) );
  OAI2BB2XL U1267 ( .B0(n1726), .B1(n1764), .A0N(\gbuff[0][7] ), .A1N(n1728), 
        .Y(n2788) );
  OAI2BB2XL U1268 ( .B0(n1726), .B1(n1763), .A0N(\gbuff[0][8] ), .A1N(n1728), 
        .Y(n2787) );
  OAI2BB2XL U1269 ( .B0(n1726), .B1(n1762), .A0N(\gbuff[0][9] ), .A1N(n1728), 
        .Y(n2786) );
  OAI2BB2XL U1270 ( .B0(n1726), .B1(n1761), .A0N(\gbuff[0][10] ), .A1N(n1728), 
        .Y(n2785) );
  OAI2BB2XL U1271 ( .B0(n1726), .B1(n1760), .A0N(\gbuff[0][11] ), .A1N(n1728), 
        .Y(n2784) );
  OAI2BB2XL U1272 ( .B0(n1726), .B1(n1759), .A0N(\gbuff[0][12] ), .A1N(n1728), 
        .Y(n2783) );
  OAI2BB2XL U1273 ( .B0(n1727), .B1(n1758), .A0N(\gbuff[0][13] ), .A1N(n1728), 
        .Y(n2782) );
  OAI2BB2XL U1274 ( .B0(n1726), .B1(n1757), .A0N(\gbuff[0][14] ), .A1N(n1728), 
        .Y(n2781) );
  OAI2BB2XL U1275 ( .B0(n1727), .B1(n1756), .A0N(\gbuff[0][15] ), .A1N(n1727), 
        .Y(n2780) );
  OAI2BB2XL U1276 ( .B0(n1726), .B1(n1755), .A0N(\gbuff[0][16] ), .A1N(n1728), 
        .Y(n2779) );
  OAI2BB2XL U1277 ( .B0(n1726), .B1(n1754), .A0N(\gbuff[0][17] ), .A1N(n1727), 
        .Y(n2778) );
  OAI2BB2XL U1278 ( .B0(n1), .B1(n1753), .A0N(\gbuff[0][18] ), .A1N(n1727), 
        .Y(n2777) );
  OAI2BB2XL U1279 ( .B0(n1726), .B1(n1752), .A0N(\gbuff[0][19] ), .A1N(n1727), 
        .Y(n2776) );
  OAI2BB2XL U1280 ( .B0(n1727), .B1(n1751), .A0N(\gbuff[0][20] ), .A1N(n1727), 
        .Y(n2775) );
  OAI2BB2XL U1281 ( .B0(n1726), .B1(n1750), .A0N(\gbuff[0][21] ), .A1N(n1727), 
        .Y(n2774) );
  OAI2BB2XL U1282 ( .B0(n1726), .B1(n1749), .A0N(\gbuff[0][22] ), .A1N(n1728), 
        .Y(n2773) );
  OAI2BB2XL U1283 ( .B0(n1727), .B1(n1747), .A0N(\gbuff[0][24] ), .A1N(n1728), 
        .Y(n2771) );
  OAI2BB2XL U1284 ( .B0(n1632), .B1(n1724), .A0N(\gbuff[1][0] ), .A1N(n1723), 
        .Y(n2763) );
  OAI2BB2XL U1285 ( .B0(n1630), .B1(n1723), .A0N(\gbuff[1][1] ), .A1N(n1724), 
        .Y(n2762) );
  OAI2BB2XL U1286 ( .B0(n1628), .B1(n1723), .A0N(\gbuff[1][2] ), .A1N(n1723), 
        .Y(n2761) );
  OAI2BB2XL U1287 ( .B0(n1626), .B1(n1723), .A0N(\gbuff[1][3] ), .A1N(n1725), 
        .Y(n2760) );
  OAI2BB2XL U1288 ( .B0(n1624), .B1(n1723), .A0N(\gbuff[1][4] ), .A1N(n1724), 
        .Y(n2759) );
  OAI2BB2XL U1289 ( .B0(n1622), .B1(n1723), .A0N(\gbuff[1][5] ), .A1N(n1725), 
        .Y(n2758) );
  OAI2BB2XL U1290 ( .B0(n1620), .B1(n1723), .A0N(\gbuff[1][6] ), .A1N(n1725), 
        .Y(n2757) );
  OAI2BB2XL U1291 ( .B0(n1618), .B1(n1723), .A0N(\gbuff[1][7] ), .A1N(n1725), 
        .Y(n2756) );
  OAI2BB2XL U1292 ( .B0(n1616), .B1(n1723), .A0N(\gbuff[1][8] ), .A1N(n1725), 
        .Y(n2755) );
  OAI2BB2XL U1293 ( .B0(n1614), .B1(n1723), .A0N(\gbuff[1][9] ), .A1N(n1725), 
        .Y(n2754) );
  OAI2BB2XL U1294 ( .B0(n1612), .B1(n1723), .A0N(\gbuff[1][10] ), .A1N(n1725), 
        .Y(n2753) );
  OAI2BB2XL U1295 ( .B0(n1610), .B1(n1723), .A0N(\gbuff[1][11] ), .A1N(n1725), 
        .Y(n2752) );
  OAI2BB2XL U1296 ( .B0(n1608), .B1(n1723), .A0N(\gbuff[1][12] ), .A1N(n1725), 
        .Y(n2751) );
  OAI2BB2XL U1297 ( .B0(n1606), .B1(n1724), .A0N(\gbuff[1][13] ), .A1N(n1725), 
        .Y(n2750) );
  OAI2BB2XL U1298 ( .B0(n1604), .B1(n1724), .A0N(\gbuff[1][14] ), .A1N(n1725), 
        .Y(n2749) );
  OAI2BB2XL U1299 ( .B0(n1602), .B1(n1724), .A0N(\gbuff[1][15] ), .A1N(n1725), 
        .Y(n2748) );
  OAI2BB2XL U1300 ( .B0(n1600), .B1(n1724), .A0N(\gbuff[1][16] ), .A1N(n1725), 
        .Y(n2747) );
  OAI2BB2XL U1301 ( .B0(n1598), .B1(n1724), .A0N(\gbuff[1][17] ), .A1N(n14), 
        .Y(n2746) );
  OAI2BB2XL U1302 ( .B0(n1596), .B1(n1724), .A0N(\gbuff[1][18] ), .A1N(n14), 
        .Y(n2745) );
  OAI2BB2XL U1303 ( .B0(n1594), .B1(n1724), .A0N(\gbuff[1][19] ), .A1N(n1725), 
        .Y(n2744) );
  OAI2BB2XL U1304 ( .B0(n1592), .B1(n1724), .A0N(\gbuff[1][20] ), .A1N(n1725), 
        .Y(n2743) );
  OAI2BB2XL U1305 ( .B0(n1590), .B1(n1724), .A0N(\gbuff[1][21] ), .A1N(n1723), 
        .Y(n2742) );
  OAI2BB2XL U1306 ( .B0(n1588), .B1(n1724), .A0N(\gbuff[1][22] ), .A1N(n1725), 
        .Y(n2741) );
  OAI2BB2XL U1307 ( .B0(n1584), .B1(n1724), .A0N(\gbuff[1][24] ), .A1N(n1725), 
        .Y(n2739) );
  OAI2BB2XL U1308 ( .B0(n1631), .B1(n1721), .A0N(\gbuff[2][0] ), .A1N(n1720), 
        .Y(n2731) );
  OAI2BB2XL U1309 ( .B0(n1629), .B1(n1720), .A0N(\gbuff[2][1] ), .A1N(n1721), 
        .Y(n2730) );
  OAI2BB2XL U1310 ( .B0(n1627), .B1(n1720), .A0N(\gbuff[2][2] ), .A1N(n1720), 
        .Y(n2729) );
  OAI2BB2XL U1311 ( .B0(n1625), .B1(n1720), .A0N(\gbuff[2][3] ), .A1N(n1722), 
        .Y(n2728) );
  OAI2BB2XL U1312 ( .B0(n1623), .B1(n1720), .A0N(\gbuff[2][4] ), .A1N(n1721), 
        .Y(n2727) );
  OAI2BB2XL U1313 ( .B0(n1621), .B1(n1720), .A0N(\gbuff[2][5] ), .A1N(n1722), 
        .Y(n2726) );
  OAI2BB2XL U1314 ( .B0(n1619), .B1(n1720), .A0N(\gbuff[2][6] ), .A1N(n1722), 
        .Y(n2725) );
  OAI2BB2XL U1315 ( .B0(n1617), .B1(n1720), .A0N(\gbuff[2][7] ), .A1N(n1722), 
        .Y(n2724) );
  OAI2BB2XL U1316 ( .B0(n1615), .B1(n1720), .A0N(\gbuff[2][8] ), .A1N(n1722), 
        .Y(n2723) );
  OAI2BB2XL U1317 ( .B0(n1613), .B1(n1720), .A0N(\gbuff[2][9] ), .A1N(n1722), 
        .Y(n2722) );
  OAI2BB2XL U1318 ( .B0(n1611), .B1(n1720), .A0N(\gbuff[2][10] ), .A1N(n1722), 
        .Y(n2721) );
  OAI2BB2XL U1319 ( .B0(n1609), .B1(n1720), .A0N(\gbuff[2][11] ), .A1N(n1722), 
        .Y(n2720) );
  OAI2BB2XL U1320 ( .B0(n1607), .B1(n1720), .A0N(\gbuff[2][12] ), .A1N(n1722), 
        .Y(n2719) );
  OAI2BB2XL U1321 ( .B0(n1605), .B1(n1721), .A0N(\gbuff[2][13] ), .A1N(n1722), 
        .Y(n2718) );
  OAI2BB2XL U1322 ( .B0(n1603), .B1(n1721), .A0N(\gbuff[2][14] ), .A1N(n1722), 
        .Y(n2717) );
  OAI2BB2XL U1323 ( .B0(n1601), .B1(n1721), .A0N(\gbuff[2][15] ), .A1N(n1722), 
        .Y(n2716) );
  OAI2BB2XL U1324 ( .B0(n1599), .B1(n1721), .A0N(\gbuff[2][16] ), .A1N(n1722), 
        .Y(n2715) );
  OAI2BB2XL U1325 ( .B0(n1597), .B1(n1721), .A0N(\gbuff[2][17] ), .A1N(n15), 
        .Y(n2714) );
  OAI2BB2XL U1326 ( .B0(n1595), .B1(n1721), .A0N(\gbuff[2][18] ), .A1N(n15), 
        .Y(n2713) );
  OAI2BB2XL U1327 ( .B0(n1593), .B1(n1721), .A0N(\gbuff[2][19] ), .A1N(n1722), 
        .Y(n2712) );
  OAI2BB2XL U1328 ( .B0(n1591), .B1(n1721), .A0N(\gbuff[2][20] ), .A1N(n1722), 
        .Y(n2711) );
  OAI2BB2XL U1329 ( .B0(n1589), .B1(n1721), .A0N(\gbuff[2][21] ), .A1N(n1720), 
        .Y(n2710) );
  OAI2BB2XL U1330 ( .B0(n1587), .B1(n1721), .A0N(\gbuff[2][22] ), .A1N(n1722), 
        .Y(n2709) );
  OAI2BB2XL U1331 ( .B0(n1583), .B1(n1721), .A0N(\gbuff[2][24] ), .A1N(n1722), 
        .Y(n2707) );
  OAI2BB2XL U1332 ( .B0(n1632), .B1(n1719), .A0N(\gbuff[3][0] ), .A1N(n1717), 
        .Y(n2699) );
  OAI2BB2XL U1333 ( .B0(n1630), .B1(n1718), .A0N(\gbuff[3][1] ), .A1N(n1717), 
        .Y(n2698) );
  OAI2BB2XL U1334 ( .B0(n1628), .B1(n1718), .A0N(\gbuff[3][2] ), .A1N(n1717), 
        .Y(n2697) );
  OAI2BB2XL U1335 ( .B0(n1626), .B1(n1718), .A0N(\gbuff[3][3] ), .A1N(n1717), 
        .Y(n2696) );
  OAI2BB2XL U1336 ( .B0(n1624), .B1(n1718), .A0N(\gbuff[3][4] ), .A1N(n1717), 
        .Y(n2695) );
  OAI2BB2XL U1337 ( .B0(n1622), .B1(n1718), .A0N(\gbuff[3][5] ), .A1N(n1717), 
        .Y(n2694) );
  OAI2BB2XL U1338 ( .B0(n1620), .B1(n1718), .A0N(\gbuff[3][6] ), .A1N(n1717), 
        .Y(n2693) );
  OAI2BB2XL U1339 ( .B0(n1618), .B1(n1718), .A0N(\gbuff[3][7] ), .A1N(n1717), 
        .Y(n2692) );
  OAI2BB2XL U1340 ( .B0(n1616), .B1(n1718), .A0N(\gbuff[3][8] ), .A1N(n1718), 
        .Y(n2691) );
  OAI2BB2XL U1341 ( .B0(n1614), .B1(n1718), .A0N(\gbuff[3][9] ), .A1N(n1719), 
        .Y(n2690) );
  OAI2BB2XL U1342 ( .B0(n1612), .B1(n1718), .A0N(\gbuff[3][10] ), .A1N(n1718), 
        .Y(n2689) );
  OAI2BB2XL U1343 ( .B0(n1610), .B1(n1718), .A0N(\gbuff[3][11] ), .A1N(n1719), 
        .Y(n2688) );
  OAI2BB2XL U1344 ( .B0(n1608), .B1(n1718), .A0N(\gbuff[3][12] ), .A1N(n1718), 
        .Y(n2687) );
  OAI2BB2XL U1345 ( .B0(n1606), .B1(n1719), .A0N(\gbuff[3][13] ), .A1N(n1719), 
        .Y(n2686) );
  OAI2BB2XL U1346 ( .B0(n1604), .B1(n1719), .A0N(\gbuff[3][14] ), .A1N(n1718), 
        .Y(n2685) );
  OAI2BB2XL U1347 ( .B0(n1602), .B1(n1719), .A0N(\gbuff[3][15] ), .A1N(n2), 
        .Y(n2684) );
  OAI2BB2XL U1348 ( .B0(n1600), .B1(n1719), .A0N(\gbuff[3][16] ), .A1N(n1719), 
        .Y(n2683) );
  OAI2BB2XL U1349 ( .B0(n1598), .B1(n1719), .A0N(\gbuff[3][17] ), .A1N(n1717), 
        .Y(n2682) );
  OAI2BB2XL U1350 ( .B0(n1596), .B1(n1719), .A0N(\gbuff[3][18] ), .A1N(n1717), 
        .Y(n2681) );
  OAI2BB2XL U1351 ( .B0(n1594), .B1(n1719), .A0N(\gbuff[3][19] ), .A1N(n1717), 
        .Y(n2680) );
  OAI2BB2XL U1352 ( .B0(n1592), .B1(n1719), .A0N(\gbuff[3][20] ), .A1N(n1717), 
        .Y(n2679) );
  OAI2BB2XL U1353 ( .B0(n1590), .B1(n1719), .A0N(\gbuff[3][21] ), .A1N(n1717), 
        .Y(n2678) );
  OAI2BB2XL U1354 ( .B0(n1588), .B1(n1719), .A0N(\gbuff[3][22] ), .A1N(n1718), 
        .Y(n2677) );
  OAI2BB2XL U1355 ( .B0(n1584), .B1(n1719), .A0N(\gbuff[3][24] ), .A1N(n1719), 
        .Y(n2675) );
  OAI2BB2XL U1356 ( .B0(n1631), .B1(n1715), .A0N(\gbuff[4][0] ), .A1N(n1714), 
        .Y(n2667) );
  OAI2BB2XL U1357 ( .B0(n1629), .B1(n1714), .A0N(\gbuff[4][1] ), .A1N(n1715), 
        .Y(n2666) );
  OAI2BB2XL U1358 ( .B0(n1627), .B1(n1714), .A0N(\gbuff[4][2] ), .A1N(n1714), 
        .Y(n2665) );
  OAI2BB2XL U1359 ( .B0(n1625), .B1(n1714), .A0N(\gbuff[4][3] ), .A1N(n1716), 
        .Y(n2664) );
  OAI2BB2XL U1360 ( .B0(n1623), .B1(n1714), .A0N(\gbuff[4][4] ), .A1N(n1715), 
        .Y(n2663) );
  OAI2BB2XL U1361 ( .B0(n1621), .B1(n1714), .A0N(\gbuff[4][5] ), .A1N(n1716), 
        .Y(n2662) );
  OAI2BB2XL U1362 ( .B0(n1619), .B1(n1714), .A0N(\gbuff[4][6] ), .A1N(n1716), 
        .Y(n2661) );
  OAI2BB2XL U1363 ( .B0(n1617), .B1(n1714), .A0N(\gbuff[4][7] ), .A1N(n1716), 
        .Y(n2660) );
  OAI2BB2XL U1364 ( .B0(n1615), .B1(n1714), .A0N(\gbuff[4][8] ), .A1N(n1716), 
        .Y(n2659) );
  OAI2BB2XL U1365 ( .B0(n1613), .B1(n1714), .A0N(\gbuff[4][9] ), .A1N(n1716), 
        .Y(n2658) );
  OAI2BB2XL U1366 ( .B0(n1611), .B1(n1714), .A0N(\gbuff[4][10] ), .A1N(n1716), 
        .Y(n2657) );
  OAI2BB2XL U1367 ( .B0(n1609), .B1(n1714), .A0N(\gbuff[4][11] ), .A1N(n1716), 
        .Y(n2656) );
  OAI2BB2XL U1368 ( .B0(n1607), .B1(n1714), .A0N(\gbuff[4][12] ), .A1N(n1716), 
        .Y(n2655) );
  OAI2BB2XL U1369 ( .B0(n1605), .B1(n1715), .A0N(\gbuff[4][13] ), .A1N(n1716), 
        .Y(n2654) );
  OAI2BB2XL U1370 ( .B0(n1603), .B1(n1715), .A0N(\gbuff[4][14] ), .A1N(n1716), 
        .Y(n2653) );
  OAI2BB2XL U1371 ( .B0(n1601), .B1(n1715), .A0N(\gbuff[4][15] ), .A1N(n1716), 
        .Y(n2652) );
  OAI2BB2XL U1372 ( .B0(n1599), .B1(n1715), .A0N(\gbuff[4][16] ), .A1N(n1716), 
        .Y(n2651) );
  OAI2BB2XL U1373 ( .B0(n1597), .B1(n1715), .A0N(\gbuff[4][17] ), .A1N(n1716), 
        .Y(n2650) );
  OAI2BB2XL U1374 ( .B0(n1595), .B1(n1715), .A0N(\gbuff[4][18] ), .A1N(n1716), 
        .Y(n2649) );
  OAI2BB2XL U1375 ( .B0(n1593), .B1(n1715), .A0N(\gbuff[4][19] ), .A1N(n16), 
        .Y(n2648) );
  OAI2BB2XL U1376 ( .B0(n1591), .B1(n1715), .A0N(\gbuff[4][20] ), .A1N(n16), 
        .Y(n2647) );
  OAI2BB2XL U1377 ( .B0(n1589), .B1(n1715), .A0N(\gbuff[4][21] ), .A1N(n16), 
        .Y(n2646) );
  OAI2BB2XL U1378 ( .B0(n1587), .B1(n1715), .A0N(\gbuff[4][22] ), .A1N(n1716), 
        .Y(n2645) );
  OAI2BB2XL U1379 ( .B0(n1583), .B1(n1715), .A0N(\gbuff[4][24] ), .A1N(n1716), 
        .Y(n2643) );
  OAI2BB2XL U1380 ( .B0(n1771), .B1(n1713), .A0N(\gbuff[5][0] ), .A1N(n1711), 
        .Y(n2635) );
  OAI2BB2XL U1381 ( .B0(n1770), .B1(n1712), .A0N(\gbuff[5][1] ), .A1N(n1711), 
        .Y(n2634) );
  OAI2BB2XL U1382 ( .B0(n1769), .B1(n1712), .A0N(\gbuff[5][2] ), .A1N(n1711), 
        .Y(n2633) );
  OAI2BB2XL U1383 ( .B0(n1768), .B1(n1712), .A0N(\gbuff[5][3] ), .A1N(n1711), 
        .Y(n2632) );
  OAI2BB2XL U1384 ( .B0(n1767), .B1(n1712), .A0N(\gbuff[5][4] ), .A1N(n1711), 
        .Y(n2631) );
  OAI2BB2XL U1385 ( .B0(n1766), .B1(n1712), .A0N(\gbuff[5][5] ), .A1N(n1711), 
        .Y(n2630) );
  OAI2BB2XL U1386 ( .B0(n1765), .B1(n1712), .A0N(\gbuff[5][6] ), .A1N(n1711), 
        .Y(n2629) );
  OAI2BB2XL U1387 ( .B0(n1764), .B1(n1712), .A0N(\gbuff[5][7] ), .A1N(n1711), 
        .Y(n2628) );
  OAI2BB2XL U1388 ( .B0(n1763), .B1(n1712), .A0N(\gbuff[5][8] ), .A1N(n1712), 
        .Y(n2627) );
  OAI2BB2XL U1389 ( .B0(n1762), .B1(n1712), .A0N(\gbuff[5][9] ), .A1N(n1713), 
        .Y(n2626) );
  OAI2BB2XL U1390 ( .B0(n1761), .B1(n1712), .A0N(\gbuff[5][10] ), .A1N(n1712), 
        .Y(n2625) );
  OAI2BB2XL U1391 ( .B0(n1760), .B1(n1712), .A0N(\gbuff[5][11] ), .A1N(n1713), 
        .Y(n2624) );
  OAI2BB2XL U1392 ( .B0(n1759), .B1(n1712), .A0N(\gbuff[5][12] ), .A1N(n1712), 
        .Y(n2623) );
  OAI2BB2XL U1393 ( .B0(n1758), .B1(n1713), .A0N(\gbuff[5][13] ), .A1N(n1713), 
        .Y(n2622) );
  OAI2BB2XL U1394 ( .B0(n1757), .B1(n1713), .A0N(\gbuff[5][14] ), .A1N(n1712), 
        .Y(n2621) );
  OAI2BB2XL U1395 ( .B0(n1756), .B1(n1713), .A0N(\gbuff[5][15] ), .A1N(n3), 
        .Y(n2620) );
  OAI2BB2XL U1396 ( .B0(n1755), .B1(n1713), .A0N(\gbuff[5][16] ), .A1N(n1713), 
        .Y(n2619) );
  OAI2BB2XL U1397 ( .B0(n1754), .B1(n1713), .A0N(\gbuff[5][17] ), .A1N(n1711), 
        .Y(n2618) );
  OAI2BB2XL U1398 ( .B0(n1753), .B1(n1713), .A0N(\gbuff[5][18] ), .A1N(n1711), 
        .Y(n2617) );
  OAI2BB2XL U1399 ( .B0(n1752), .B1(n1713), .A0N(\gbuff[5][19] ), .A1N(n1711), 
        .Y(n2616) );
  OAI2BB2XL U1400 ( .B0(n1751), .B1(n1713), .A0N(\gbuff[5][20] ), .A1N(n1711), 
        .Y(n2615) );
  OAI2BB2XL U1401 ( .B0(n1750), .B1(n1713), .A0N(\gbuff[5][21] ), .A1N(n1711), 
        .Y(n2614) );
  OAI2BB2XL U1402 ( .B0(n1749), .B1(n1713), .A0N(\gbuff[5][22] ), .A1N(n1712), 
        .Y(n2613) );
  OAI2BB2XL U1403 ( .B0(n1747), .B1(n1713), .A0N(\gbuff[5][24] ), .A1N(n1713), 
        .Y(n2611) );
  OAI2BB2XL U1404 ( .B0(n1771), .B1(n1710), .A0N(\gbuff[6][0] ), .A1N(n1708), 
        .Y(n2603) );
  OAI2BB2XL U1405 ( .B0(n1770), .B1(n1709), .A0N(\gbuff[6][1] ), .A1N(n1708), 
        .Y(n2602) );
  OAI2BB2XL U1406 ( .B0(n1769), .B1(n1709), .A0N(\gbuff[6][2] ), .A1N(n1708), 
        .Y(n2601) );
  OAI2BB2XL U1407 ( .B0(n1768), .B1(n1709), .A0N(\gbuff[6][3] ), .A1N(n1708), 
        .Y(n2600) );
  OAI2BB2XL U1408 ( .B0(n1767), .B1(n1709), .A0N(\gbuff[6][4] ), .A1N(n1708), 
        .Y(n2599) );
  OAI2BB2XL U1409 ( .B0(n1766), .B1(n1709), .A0N(\gbuff[6][5] ), .A1N(n1708), 
        .Y(n2598) );
  OAI2BB2XL U1410 ( .B0(n1765), .B1(n1709), .A0N(\gbuff[6][6] ), .A1N(n1708), 
        .Y(n2597) );
  OAI2BB2XL U1411 ( .B0(n1764), .B1(n1709), .A0N(\gbuff[6][7] ), .A1N(n1708), 
        .Y(n2596) );
  OAI2BB2XL U1412 ( .B0(n1763), .B1(n1709), .A0N(\gbuff[6][8] ), .A1N(n1709), 
        .Y(n2595) );
  OAI2BB2XL U1413 ( .B0(n1762), .B1(n1709), .A0N(\gbuff[6][9] ), .A1N(n1710), 
        .Y(n2594) );
  OAI2BB2XL U1414 ( .B0(n1761), .B1(n1709), .A0N(\gbuff[6][10] ), .A1N(n1709), 
        .Y(n2593) );
  OAI2BB2XL U1415 ( .B0(n1760), .B1(n1709), .A0N(\gbuff[6][11] ), .A1N(n1710), 
        .Y(n2592) );
  OAI2BB2XL U1416 ( .B0(n1759), .B1(n1709), .A0N(\gbuff[6][12] ), .A1N(n1709), 
        .Y(n2591) );
  OAI2BB2XL U1417 ( .B0(n1758), .B1(n1710), .A0N(\gbuff[6][13] ), .A1N(n1710), 
        .Y(n2590) );
  OAI2BB2XL U1418 ( .B0(n1757), .B1(n1710), .A0N(\gbuff[6][14] ), .A1N(n1709), 
        .Y(n2589) );
  OAI2BB2XL U1419 ( .B0(n1756), .B1(n1710), .A0N(\gbuff[6][15] ), .A1N(n4), 
        .Y(n2588) );
  OAI2BB2XL U1420 ( .B0(n1755), .B1(n1710), .A0N(\gbuff[6][16] ), .A1N(n1710), 
        .Y(n2587) );
  OAI2BB2XL U1421 ( .B0(n1754), .B1(n1710), .A0N(\gbuff[6][17] ), .A1N(n1708), 
        .Y(n2586) );
  OAI2BB2XL U1422 ( .B0(n1753), .B1(n1710), .A0N(\gbuff[6][18] ), .A1N(n1708), 
        .Y(n2585) );
  OAI2BB2XL U1423 ( .B0(n1752), .B1(n1710), .A0N(\gbuff[6][19] ), .A1N(n1708), 
        .Y(n2584) );
  OAI2BB2XL U1424 ( .B0(n1751), .B1(n1710), .A0N(\gbuff[6][20] ), .A1N(n1708), 
        .Y(n2583) );
  OAI2BB2XL U1425 ( .B0(n1750), .B1(n1710), .A0N(\gbuff[6][21] ), .A1N(n1708), 
        .Y(n2582) );
  OAI2BB2XL U1426 ( .B0(n1749), .B1(n1710), .A0N(\gbuff[6][22] ), .A1N(n1709), 
        .Y(n2581) );
  OAI2BB2XL U1427 ( .B0(n1747), .B1(n1710), .A0N(\gbuff[6][24] ), .A1N(n1710), 
        .Y(n2579) );
  OAI2BB2XL U1428 ( .B0(n1771), .B1(n1707), .A0N(\gbuff[7][0] ), .A1N(n1705), 
        .Y(n2571) );
  OAI2BB2XL U1429 ( .B0(n1770), .B1(n1706), .A0N(\gbuff[7][1] ), .A1N(n1705), 
        .Y(n2570) );
  OAI2BB2XL U1430 ( .B0(n1769), .B1(n1706), .A0N(\gbuff[7][2] ), .A1N(n1705), 
        .Y(n2569) );
  OAI2BB2XL U1431 ( .B0(n1768), .B1(n1706), .A0N(\gbuff[7][3] ), .A1N(n1705), 
        .Y(n2568) );
  OAI2BB2XL U1432 ( .B0(n1767), .B1(n1706), .A0N(\gbuff[7][4] ), .A1N(n1705), 
        .Y(n2567) );
  OAI2BB2XL U1433 ( .B0(n1766), .B1(n1706), .A0N(\gbuff[7][5] ), .A1N(n1705), 
        .Y(n2566) );
  OAI2BB2XL U1434 ( .B0(n1765), .B1(n1706), .A0N(\gbuff[7][6] ), .A1N(n1705), 
        .Y(n2565) );
  OAI2BB2XL U1435 ( .B0(n1764), .B1(n1706), .A0N(\gbuff[7][7] ), .A1N(n1705), 
        .Y(n2564) );
  OAI2BB2XL U1436 ( .B0(n1763), .B1(n1706), .A0N(\gbuff[7][8] ), .A1N(n1706), 
        .Y(n2563) );
  OAI2BB2XL U1437 ( .B0(n1762), .B1(n1706), .A0N(\gbuff[7][9] ), .A1N(n1707), 
        .Y(n2562) );
  OAI2BB2XL U1438 ( .B0(n1761), .B1(n1706), .A0N(\gbuff[7][10] ), .A1N(n1706), 
        .Y(n2561) );
  OAI2BB2XL U1439 ( .B0(n1760), .B1(n1706), .A0N(\gbuff[7][11] ), .A1N(n1707), 
        .Y(n2560) );
  OAI2BB2XL U1440 ( .B0(n1759), .B1(n1706), .A0N(\gbuff[7][12] ), .A1N(n1706), 
        .Y(n2559) );
  OAI2BB2XL U1441 ( .B0(n1758), .B1(n1707), .A0N(\gbuff[7][13] ), .A1N(n1707), 
        .Y(n2558) );
  OAI2BB2XL U1442 ( .B0(n1757), .B1(n1707), .A0N(\gbuff[7][14] ), .A1N(n1706), 
        .Y(n2557) );
  OAI2BB2XL U1443 ( .B0(n1756), .B1(n1707), .A0N(\gbuff[7][15] ), .A1N(n5), 
        .Y(n2556) );
  OAI2BB2XL U1444 ( .B0(n1755), .B1(n1707), .A0N(\gbuff[7][16] ), .A1N(n1707), 
        .Y(n2555) );
  OAI2BB2XL U1445 ( .B0(n1754), .B1(n1707), .A0N(\gbuff[7][17] ), .A1N(n1705), 
        .Y(n2554) );
  OAI2BB2XL U1446 ( .B0(n1753), .B1(n1707), .A0N(\gbuff[7][18] ), .A1N(n1705), 
        .Y(n2553) );
  OAI2BB2XL U1447 ( .B0(n1752), .B1(n1707), .A0N(\gbuff[7][19] ), .A1N(n1705), 
        .Y(n2552) );
  OAI2BB2XL U1448 ( .B0(n1751), .B1(n1707), .A0N(\gbuff[7][20] ), .A1N(n1705), 
        .Y(n2551) );
  OAI2BB2XL U1449 ( .B0(n1750), .B1(n1707), .A0N(\gbuff[7][21] ), .A1N(n1705), 
        .Y(n2550) );
  OAI2BB2XL U1450 ( .B0(n1749), .B1(n1707), .A0N(\gbuff[7][22] ), .A1N(n1706), 
        .Y(n2549) );
  OAI2BB2XL U1451 ( .B0(n1747), .B1(n1707), .A0N(\gbuff[7][24] ), .A1N(n1707), 
        .Y(n2547) );
  MX4X1 U1452 ( .A(\gbuff[4][0] ), .B(\gbuff[5][0] ), .C(\gbuff[6][0] ), .D(
        \gbuff[7][0] ), .S0(n1436), .S1(n1398), .Y(n23) );
  MX4X1 U1453 ( .A(\gbuff[20][0] ), .B(\gbuff[21][0] ), .C(\gbuff[22][0] ), 
        .D(\gbuff[23][0] ), .S0(n1437), .S1(n1398), .Y(n19) );
  MX4X1 U1454 ( .A(\gbuff[4][1] ), .B(\gbuff[5][1] ), .C(\gbuff[6][1] ), .D(
        \gbuff[7][1] ), .S0(n1418), .S1(n1399), .Y(n33) );
  MX4X1 U1455 ( .A(\gbuff[20][1] ), .B(\gbuff[21][1] ), .C(\gbuff[22][1] ), 
        .D(\gbuff[23][1] ), .S0(n1418), .S1(n1399), .Y(n29) );
  MX4X1 U1456 ( .A(\gbuff[4][2] ), .B(\gbuff[5][2] ), .C(\gbuff[6][2] ), .D(
        \gbuff[7][2] ), .S0(n1419), .S1(n1400), .Y(n43) );
  MX4X1 U1457 ( .A(\gbuff[20][2] ), .B(\gbuff[21][2] ), .C(\gbuff[22][2] ), 
        .D(\gbuff[23][2] ), .S0(n1418), .S1(n1399), .Y(n39) );
  MX4X1 U1458 ( .A(\gbuff[4][3] ), .B(\gbuff[5][3] ), .C(\gbuff[6][3] ), .D(
        \gbuff[7][3] ), .S0(n1419), .S1(n1400), .Y(n53) );
  MX4X1 U1459 ( .A(\gbuff[20][3] ), .B(\gbuff[21][3] ), .C(\gbuff[22][3] ), 
        .D(\gbuff[23][3] ), .S0(n1419), .S1(n1400), .Y(n49) );
  MX4X1 U1460 ( .A(\gbuff[4][4] ), .B(\gbuff[5][4] ), .C(\gbuff[6][4] ), .D(
        \gbuff[7][4] ), .S0(n1420), .S1(n1401), .Y(n63) );
  MX4X1 U1461 ( .A(\gbuff[20][4] ), .B(\gbuff[21][4] ), .C(\gbuff[22][4] ), 
        .D(\gbuff[23][4] ), .S0(n1419), .S1(n1400), .Y(n59) );
  MX4X1 U1462 ( .A(\gbuff[4][5] ), .B(\gbuff[5][5] ), .C(\gbuff[6][5] ), .D(
        \gbuff[7][5] ), .S0(n1420), .S1(n1401), .Y(n73) );
  MX4X1 U1463 ( .A(\gbuff[20][5] ), .B(\gbuff[21][5] ), .C(\gbuff[22][5] ), 
        .D(\gbuff[23][5] ), .S0(n1420), .S1(n1401), .Y(n69) );
  MX4X1 U1464 ( .A(\gbuff[4][6] ), .B(\gbuff[5][6] ), .C(\gbuff[6][6] ), .D(
        \gbuff[7][6] ), .S0(n1421), .S1(n1402), .Y(n83) );
  MX4X1 U1465 ( .A(\gbuff[20][6] ), .B(\gbuff[21][6] ), .C(\gbuff[22][6] ), 
        .D(\gbuff[23][6] ), .S0(n1421), .S1(n1402), .Y(n79) );
  MX4X1 U1466 ( .A(\gbuff[4][7] ), .B(\gbuff[5][7] ), .C(\gbuff[6][7] ), .D(
        \gbuff[7][7] ), .S0(n1436), .S1(n1403), .Y(n93) );
  MX4X1 U1467 ( .A(\gbuff[20][7] ), .B(\gbuff[21][7] ), .C(\gbuff[22][7] ), 
        .D(\gbuff[23][7] ), .S0(n1421), .S1(n1402), .Y(n89) );
  MX4X1 U1468 ( .A(\gbuff[4][8] ), .B(\gbuff[5][8] ), .C(\gbuff[6][8] ), .D(
        \gbuff[7][8] ), .S0(n1436), .S1(n1403), .Y(n106) );
  MX4X1 U1469 ( .A(\gbuff[20][8] ), .B(\gbuff[21][8] ), .C(\gbuff[22][8] ), 
        .D(\gbuff[23][8] ), .S0(n1437), .S1(n1403), .Y(n99) );
  MX4X1 U1470 ( .A(\gbuff[4][9] ), .B(\gbuff[5][9] ), .C(\gbuff[6][9] ), .D(
        \gbuff[7][9] ), .S0(n1422), .S1(n1404), .Y(n124) );
  MX4X1 U1471 ( .A(\gbuff[20][9] ), .B(\gbuff[21][9] ), .C(\gbuff[22][9] ), 
        .D(\gbuff[23][9] ), .S0(n1422), .S1(n1404), .Y(n119) );
  MX4X1 U1472 ( .A(\gbuff[4][10] ), .B(\gbuff[5][10] ), .C(\gbuff[6][10] ), 
        .D(\gbuff[7][10] ), .S0(n1422), .S1(n1404), .Y(n1176) );
  MX4X1 U1473 ( .A(\gbuff[20][10] ), .B(\gbuff[21][10] ), .C(\gbuff[22][10] ), 
        .D(\gbuff[23][10] ), .S0(n1422), .S1(n1404), .Y(n1172) );
  MX4X1 U1474 ( .A(\gbuff[4][11] ), .B(\gbuff[5][11] ), .C(\gbuff[6][11] ), 
        .D(\gbuff[7][11] ), .S0(n1423), .S1(n1405), .Y(n1186) );
  MX4X1 U1475 ( .A(\gbuff[20][11] ), .B(\gbuff[21][11] ), .C(\gbuff[22][11] ), 
        .D(\gbuff[23][11] ), .S0(n1423), .S1(n1405), .Y(n1182) );
  MX4X1 U1476 ( .A(\gbuff[4][12] ), .B(\gbuff[5][12] ), .C(\gbuff[6][12] ), 
        .D(\gbuff[7][12] ), .S0(n1424), .S1(n1406), .Y(n1196) );
  MX4X1 U1477 ( .A(\gbuff[20][12] ), .B(\gbuff[21][12] ), .C(\gbuff[22][12] ), 
        .D(\gbuff[23][12] ), .S0(n1423), .S1(n1405), .Y(n1192) );
  MX4X1 U1478 ( .A(\gbuff[4][13] ), .B(\gbuff[5][13] ), .C(\gbuff[6][13] ), 
        .D(\gbuff[7][13] ), .S0(n1424), .S1(n1406), .Y(n1206) );
  MX4X1 U1479 ( .A(\gbuff[20][13] ), .B(\gbuff[21][13] ), .C(\gbuff[22][13] ), 
        .D(\gbuff[23][13] ), .S0(n1424), .S1(n1406), .Y(n1202) );
  MX4X1 U1480 ( .A(\gbuff[4][14] ), .B(\gbuff[5][14] ), .C(\gbuff[6][14] ), 
        .D(\gbuff[7][14] ), .S0(n1425), .S1(n1407), .Y(n1216) );
  MX4X1 U1481 ( .A(\gbuff[20][14] ), .B(\gbuff[21][14] ), .C(\gbuff[22][14] ), 
        .D(\gbuff[23][14] ), .S0(n1425), .S1(n1407), .Y(n1212) );
  MX4X1 U1482 ( .A(\gbuff[4][15] ), .B(\gbuff[5][15] ), .C(\gbuff[6][15] ), 
        .D(\gbuff[7][15] ), .S0(n1426), .S1(n1408), .Y(n1226) );
  MX4X1 U1483 ( .A(\gbuff[20][15] ), .B(\gbuff[21][15] ), .C(\gbuff[22][15] ), 
        .D(\gbuff[23][15] ), .S0(n1425), .S1(n1407), .Y(n1222) );
  MX4X1 U1484 ( .A(\gbuff[4][16] ), .B(\gbuff[5][16] ), .C(\gbuff[6][16] ), 
        .D(\gbuff[7][16] ), .S0(n1426), .S1(n1408), .Y(n1236) );
  MX4X1 U1485 ( .A(\gbuff[20][16] ), .B(\gbuff[21][16] ), .C(\gbuff[22][16] ), 
        .D(\gbuff[23][16] ), .S0(n1426), .S1(n1408), .Y(n1232) );
  MX4X1 U1486 ( .A(\gbuff[4][17] ), .B(\gbuff[5][17] ), .C(\gbuff[6][17] ), 
        .D(\gbuff[7][17] ), .S0(n1427), .S1(n1409), .Y(n1246) );
  MX4X1 U1487 ( .A(\gbuff[20][17] ), .B(\gbuff[21][17] ), .C(\gbuff[22][17] ), 
        .D(\gbuff[23][17] ), .S0(n1426), .S1(n1408), .Y(n1242) );
  MX4X1 U1488 ( .A(\gbuff[4][18] ), .B(\gbuff[5][18] ), .C(\gbuff[6][18] ), 
        .D(\gbuff[7][18] ), .S0(n1427), .S1(n1409), .Y(n1256) );
  MX4X1 U1489 ( .A(\gbuff[20][18] ), .B(\gbuff[21][18] ), .C(\gbuff[22][18] ), 
        .D(\gbuff[23][18] ), .S0(n1427), .S1(n1409), .Y(n1252) );
  MX4X1 U1490 ( .A(\gbuff[4][19] ), .B(\gbuff[5][19] ), .C(\gbuff[6][19] ), 
        .D(\gbuff[7][19] ), .S0(n1428), .S1(n1410), .Y(n1266) );
  MX4X1 U1491 ( .A(\gbuff[20][19] ), .B(\gbuff[21][19] ), .C(\gbuff[22][19] ), 
        .D(\gbuff[23][19] ), .S0(n1428), .S1(n1410), .Y(n1262) );
  MX4X1 U1492 ( .A(\gbuff[4][20] ), .B(\gbuff[5][20] ), .C(\gbuff[6][20] ), 
        .D(\gbuff[7][20] ), .S0(n1429), .S1(n1411), .Y(n1276) );
  MX4X1 U1493 ( .A(\gbuff[20][20] ), .B(\gbuff[21][20] ), .C(\gbuff[22][20] ), 
        .D(\gbuff[23][20] ), .S0(n1428), .S1(n1410), .Y(n1272) );
  MX4X1 U1494 ( .A(\gbuff[4][21] ), .B(\gbuff[5][21] ), .C(\gbuff[6][21] ), 
        .D(\gbuff[7][21] ), .S0(n1429), .S1(n1411), .Y(n1286) );
  MX4X1 U1495 ( .A(\gbuff[20][21] ), .B(\gbuff[21][21] ), .C(\gbuff[22][21] ), 
        .D(\gbuff[23][21] ), .S0(n1429), .S1(n1411), .Y(n1282) );
  MX4X1 U1496 ( .A(\gbuff[4][22] ), .B(\gbuff[5][22] ), .C(\gbuff[6][22] ), 
        .D(\gbuff[7][22] ), .S0(n1430), .S1(n1412), .Y(n1296) );
  MX4X1 U1497 ( .A(\gbuff[20][22] ), .B(\gbuff[21][22] ), .C(\gbuff[22][22] ), 
        .D(\gbuff[23][22] ), .S0(n1430), .S1(n1412), .Y(n1292) );
  MX4X1 U1498 ( .A(\gbuff[4][23] ), .B(\gbuff[5][23] ), .C(\gbuff[6][23] ), 
        .D(\gbuff[7][23] ), .S0(n1430), .S1(n1412), .Y(n1306) );
  MX4X1 U1499 ( .A(\gbuff[20][23] ), .B(\gbuff[21][23] ), .C(\gbuff[22][23] ), 
        .D(\gbuff[23][23] ), .S0(n1430), .S1(n1412), .Y(n1302) );
  MX4X1 U1500 ( .A(\gbuff[4][24] ), .B(\gbuff[5][24] ), .C(\gbuff[6][24] ), 
        .D(\gbuff[7][24] ), .S0(n1431), .S1(n1413), .Y(n1316) );
  MX4X1 U1501 ( .A(\gbuff[20][24] ), .B(\gbuff[21][24] ), .C(\gbuff[22][24] ), 
        .D(\gbuff[23][24] ), .S0(n1431), .S1(n1413), .Y(n1312) );
  MX4X1 U1502 ( .A(\gbuff[4][25] ), .B(\gbuff[5][25] ), .C(\gbuff[6][25] ), 
        .D(\gbuff[7][25] ), .S0(n1432), .S1(n1414), .Y(n1326) );
  MX4X1 U1503 ( .A(\gbuff[20][25] ), .B(\gbuff[21][25] ), .C(\gbuff[22][25] ), 
        .D(\gbuff[23][25] ), .S0(n1431), .S1(n1413), .Y(n1322) );
  MX4X1 U1504 ( .A(\gbuff[4][26] ), .B(\gbuff[5][26] ), .C(\gbuff[6][26] ), 
        .D(\gbuff[7][26] ), .S0(n1432), .S1(n1414), .Y(n1336) );
  MX4X1 U1505 ( .A(\gbuff[20][26] ), .B(\gbuff[21][26] ), .C(\gbuff[22][26] ), 
        .D(\gbuff[23][26] ), .S0(n1432), .S1(n1414), .Y(n1332) );
  MX4X1 U1506 ( .A(\gbuff[4][27] ), .B(\gbuff[5][27] ), .C(\gbuff[6][27] ), 
        .D(\gbuff[7][27] ), .S0(n1433), .S1(n1415), .Y(n1346) );
  MX4X1 U1507 ( .A(\gbuff[20][27] ), .B(\gbuff[21][27] ), .C(\gbuff[22][27] ), 
        .D(\gbuff[23][27] ), .S0(n1433), .S1(n1415), .Y(n1342) );
  MX4X1 U1508 ( .A(\gbuff[4][28] ), .B(\gbuff[5][28] ), .C(\gbuff[6][28] ), 
        .D(\gbuff[7][28] ), .S0(n1434), .S1(n1416), .Y(n1356) );
  MX4X1 U1509 ( .A(\gbuff[20][28] ), .B(\gbuff[21][28] ), .C(\gbuff[22][28] ), 
        .D(\gbuff[23][28] ), .S0(n1433), .S1(n1415), .Y(n1352) );
  MX4X1 U1510 ( .A(\gbuff[4][29] ), .B(\gbuff[5][29] ), .C(\gbuff[6][29] ), 
        .D(\gbuff[7][29] ), .S0(n1434), .S1(n1416), .Y(n1366) );
  MX4X1 U1511 ( .A(\gbuff[20][29] ), .B(\gbuff[21][29] ), .C(\gbuff[22][29] ), 
        .D(\gbuff[23][29] ), .S0(n1434), .S1(n1416), .Y(n1362) );
  MX4X1 U1512 ( .A(\gbuff[4][30] ), .B(\gbuff[5][30] ), .C(\gbuff[6][30] ), 
        .D(\gbuff[7][30] ), .S0(n1435), .S1(n1404), .Y(n1376) );
  MX4X1 U1513 ( .A(\gbuff[20][30] ), .B(\gbuff[21][30] ), .C(\gbuff[22][30] ), 
        .D(\gbuff[23][30] ), .S0(n1434), .S1(n1416), .Y(n1372) );
  MX4X1 U1514 ( .A(\gbuff[4][31] ), .B(\gbuff[5][31] ), .C(\gbuff[6][31] ), 
        .D(\gbuff[7][31] ), .S0(n1435), .S1(n1406), .Y(n1386) );
  MX4X1 U1515 ( .A(\gbuff[20][31] ), .B(\gbuff[21][31] ), .C(\gbuff[22][31] ), 
        .D(\gbuff[23][31] ), .S0(n1435), .S1(n1403), .Y(n1382) );
  MX4X1 U1516 ( .A(\gbuff[0][0] ), .B(\gbuff[1][0] ), .C(\gbuff[2][0] ), .D(
        \gbuff[3][0] ), .S0(n1436), .S1(n1398), .Y(n24) );
  MX4X1 U1517 ( .A(\gbuff[16][0] ), .B(\gbuff[17][0] ), .C(\gbuff[18][0] ), 
        .D(\gbuff[19][0] ), .S0(n1436), .S1(n1398), .Y(n20) );
  MX4X1 U1518 ( .A(\gbuff[0][1] ), .B(\gbuff[1][1] ), .C(\gbuff[2][1] ), .D(
        \gbuff[3][1] ), .S0(n1418), .S1(n1399), .Y(n34) );
  MX4X1 U1519 ( .A(\gbuff[16][1] ), .B(\gbuff[17][1] ), .C(\gbuff[18][1] ), 
        .D(\gbuff[19][1] ), .S0(n1418), .S1(n1399), .Y(n30) );
  MX4X1 U1520 ( .A(\gbuff[0][2] ), .B(\gbuff[1][2] ), .C(\gbuff[2][2] ), .D(
        \gbuff[3][2] ), .S0(n1419), .S1(n1400), .Y(n44) );
  MX4X1 U1521 ( .A(\gbuff[16][2] ), .B(\gbuff[17][2] ), .C(\gbuff[18][2] ), 
        .D(\gbuff[19][2] ), .S0(n1418), .S1(n1399), .Y(n40) );
  MX4X1 U1522 ( .A(\gbuff[0][3] ), .B(\gbuff[1][3] ), .C(\gbuff[2][3] ), .D(
        \gbuff[3][3] ), .S0(n1419), .S1(n1400), .Y(n54) );
  MX4X1 U1523 ( .A(\gbuff[16][3] ), .B(\gbuff[17][3] ), .C(\gbuff[18][3] ), 
        .D(\gbuff[19][3] ), .S0(n1419), .S1(n1400), .Y(n50) );
  MX4X1 U1524 ( .A(\gbuff[0][4] ), .B(\gbuff[1][4] ), .C(\gbuff[2][4] ), .D(
        \gbuff[3][4] ), .S0(n1420), .S1(n1401), .Y(n64) );
  MX4X1 U1525 ( .A(\gbuff[16][4] ), .B(\gbuff[17][4] ), .C(\gbuff[18][4] ), 
        .D(\gbuff[19][4] ), .S0(n1420), .S1(n1401), .Y(n60) );
  MX4X1 U1526 ( .A(\gbuff[0][5] ), .B(\gbuff[1][5] ), .C(\gbuff[2][5] ), .D(
        \gbuff[3][5] ), .S0(n1420), .S1(n1401), .Y(n74) );
  MX4X1 U1527 ( .A(\gbuff[16][5] ), .B(\gbuff[17][5] ), .C(\gbuff[18][5] ), 
        .D(\gbuff[19][5] ), .S0(n1420), .S1(n1401), .Y(n70) );
  MX4X1 U1528 ( .A(\gbuff[0][6] ), .B(\gbuff[1][6] ), .C(\gbuff[2][6] ), .D(
        \gbuff[3][6] ), .S0(n1421), .S1(n1402), .Y(n84) );
  MX4X1 U1529 ( .A(\gbuff[16][6] ), .B(\gbuff[17][6] ), .C(\gbuff[18][6] ), 
        .D(\gbuff[19][6] ), .S0(n1421), .S1(n1402), .Y(n80) );
  MX4X1 U1530 ( .A(\gbuff[0][7] ), .B(\gbuff[1][7] ), .C(\gbuff[2][7] ), .D(
        \gbuff[3][7] ), .S0(n1436), .S1(n1403), .Y(n94) );
  MX4X1 U1531 ( .A(\gbuff[16][7] ), .B(\gbuff[17][7] ), .C(\gbuff[18][7] ), 
        .D(\gbuff[19][7] ), .S0(n1421), .S1(n1402), .Y(n90) );
  MX4X1 U1532 ( .A(\gbuff[0][8] ), .B(\gbuff[1][8] ), .C(\gbuff[2][8] ), .D(
        \gbuff[3][8] ), .S0(n1436), .S1(n1403), .Y(n108) );
  MX4X1 U1533 ( .A(\gbuff[16][8] ), .B(\gbuff[17][8] ), .C(\gbuff[18][8] ), 
        .D(\gbuff[19][8] ), .S0(n1437), .S1(n1403), .Y(n100) );
  MX4X1 U1534 ( .A(\gbuff[0][9] ), .B(\gbuff[1][9] ), .C(\gbuff[2][9] ), .D(
        \gbuff[3][9] ), .S0(n1422), .S1(n1404), .Y(n125) );
  MX4X1 U1535 ( .A(\gbuff[16][9] ), .B(\gbuff[17][9] ), .C(\gbuff[18][9] ), 
        .D(\gbuff[19][9] ), .S0(n1422), .S1(n1404), .Y(n121) );
  MX4X1 U1536 ( .A(\gbuff[0][10] ), .B(\gbuff[1][10] ), .C(\gbuff[2][10] ), 
        .D(\gbuff[3][10] ), .S0(n1423), .S1(n1405), .Y(n1177) );
  MX4X1 U1537 ( .A(\gbuff[16][10] ), .B(\gbuff[17][10] ), .C(\gbuff[18][10] ), 
        .D(\gbuff[19][10] ), .S0(n1422), .S1(n1404), .Y(n1173) );
  MX4X1 U1538 ( .A(\gbuff[0][11] ), .B(\gbuff[1][11] ), .C(\gbuff[2][11] ), 
        .D(\gbuff[3][11] ), .S0(n1423), .S1(n1405), .Y(n1187) );
  MX4X1 U1539 ( .A(\gbuff[16][11] ), .B(\gbuff[17][11] ), .C(\gbuff[18][11] ), 
        .D(\gbuff[19][11] ), .S0(n1423), .S1(n1405), .Y(n1183) );
  MX4X1 U1540 ( .A(\gbuff[0][12] ), .B(\gbuff[1][12] ), .C(\gbuff[2][12] ), 
        .D(\gbuff[3][12] ), .S0(n1424), .S1(n1406), .Y(n1197) );
  MX4X1 U1541 ( .A(\gbuff[16][12] ), .B(\gbuff[17][12] ), .C(\gbuff[18][12] ), 
        .D(\gbuff[19][12] ), .S0(n1423), .S1(n1405), .Y(n1193) );
  MX4X1 U1542 ( .A(\gbuff[0][13] ), .B(\gbuff[1][13] ), .C(\gbuff[2][13] ), 
        .D(\gbuff[3][13] ), .S0(n1424), .S1(n1406), .Y(n1207) );
  MX4X1 U1543 ( .A(\gbuff[16][13] ), .B(\gbuff[17][13] ), .C(\gbuff[18][13] ), 
        .D(\gbuff[19][13] ), .S0(n1424), .S1(n1406), .Y(n1203) );
  MX4X1 U1544 ( .A(\gbuff[0][14] ), .B(\gbuff[1][14] ), .C(\gbuff[2][14] ), 
        .D(\gbuff[3][14] ), .S0(n1425), .S1(n1407), .Y(n1217) );
  MX4X1 U1545 ( .A(\gbuff[16][14] ), .B(\gbuff[17][14] ), .C(\gbuff[18][14] ), 
        .D(\gbuff[19][14] ), .S0(n1425), .S1(n1407), .Y(n1213) );
  MX4X1 U1546 ( .A(\gbuff[0][15] ), .B(\gbuff[1][15] ), .C(\gbuff[2][15] ), 
        .D(\gbuff[3][15] ), .S0(n1426), .S1(n1408), .Y(n1227) );
  MX4X1 U1547 ( .A(\gbuff[16][15] ), .B(\gbuff[17][15] ), .C(\gbuff[18][15] ), 
        .D(\gbuff[19][15] ), .S0(n1425), .S1(n1407), .Y(n1223) );
  MX4X1 U1548 ( .A(\gbuff[0][16] ), .B(\gbuff[1][16] ), .C(\gbuff[2][16] ), 
        .D(\gbuff[3][16] ), .S0(n1426), .S1(n1408), .Y(n1237) );
  MX4X1 U1549 ( .A(\gbuff[16][16] ), .B(\gbuff[17][16] ), .C(\gbuff[18][16] ), 
        .D(\gbuff[19][16] ), .S0(n1426), .S1(n1408), .Y(n1233) );
  MX4X1 U1550 ( .A(\gbuff[0][17] ), .B(\gbuff[1][17] ), .C(\gbuff[2][17] ), 
        .D(\gbuff[3][17] ), .S0(n1427), .S1(n1409), .Y(n1247) );
  MX4X1 U1551 ( .A(\gbuff[16][17] ), .B(\gbuff[17][17] ), .C(\gbuff[18][17] ), 
        .D(\gbuff[19][17] ), .S0(n1427), .S1(n1409), .Y(n1243) );
  MX4X1 U1552 ( .A(\gbuff[0][18] ), .B(\gbuff[1][18] ), .C(\gbuff[2][18] ), 
        .D(\gbuff[3][18] ), .S0(n1427), .S1(n1409), .Y(n1257) );
  MX4X1 U1553 ( .A(\gbuff[16][18] ), .B(\gbuff[17][18] ), .C(\gbuff[18][18] ), 
        .D(\gbuff[19][18] ), .S0(n1427), .S1(n1409), .Y(n1253) );
  MX4X1 U1554 ( .A(\gbuff[0][19] ), .B(\gbuff[1][19] ), .C(\gbuff[2][19] ), 
        .D(\gbuff[3][19] ), .S0(n1428), .S1(n1410), .Y(n1267) );
  MX4X1 U1555 ( .A(\gbuff[16][19] ), .B(\gbuff[17][19] ), .C(\gbuff[18][19] ), 
        .D(\gbuff[19][19] ), .S0(n1428), .S1(n1410), .Y(n1263) );
  MX4X1 U1556 ( .A(\gbuff[0][20] ), .B(\gbuff[1][20] ), .C(\gbuff[2][20] ), 
        .D(\gbuff[3][20] ), .S0(n1429), .S1(n1411), .Y(n1277) );
  MX4X1 U1557 ( .A(\gbuff[16][20] ), .B(\gbuff[17][20] ), .C(\gbuff[18][20] ), 
        .D(\gbuff[19][20] ), .S0(n1428), .S1(n1410), .Y(n1273) );
  MX4X1 U1558 ( .A(\gbuff[0][21] ), .B(\gbuff[1][21] ), .C(\gbuff[2][21] ), 
        .D(\gbuff[3][21] ), .S0(n1429), .S1(n1411), .Y(n1287) );
  MX4X1 U1559 ( .A(\gbuff[16][21] ), .B(\gbuff[17][21] ), .C(\gbuff[18][21] ), 
        .D(\gbuff[19][21] ), .S0(n1429), .S1(n1411), .Y(n1283) );
  MX4X1 U1560 ( .A(\gbuff[0][22] ), .B(\gbuff[1][22] ), .C(\gbuff[2][22] ), 
        .D(\gbuff[3][22] ), .S0(n1430), .S1(n1412), .Y(n1297) );
  MX4X1 U1561 ( .A(\gbuff[16][22] ), .B(\gbuff[17][22] ), .C(\gbuff[18][22] ), 
        .D(\gbuff[19][22] ), .S0(n1430), .S1(n1412), .Y(n1293) );
  MX4X1 U1562 ( .A(\gbuff[0][23] ), .B(\gbuff[1][23] ), .C(\gbuff[2][23] ), 
        .D(\gbuff[3][23] ), .S0(n1431), .S1(n1413), .Y(n1307) );
  MX4X1 U1563 ( .A(\gbuff[16][23] ), .B(\gbuff[17][23] ), .C(\gbuff[18][23] ), 
        .D(\gbuff[19][23] ), .S0(n1430), .S1(n1412), .Y(n1303) );
  MX4X1 U1564 ( .A(\gbuff[0][24] ), .B(\gbuff[1][24] ), .C(\gbuff[2][24] ), 
        .D(\gbuff[3][24] ), .S0(n1431), .S1(n1413), .Y(n1317) );
  MX4X1 U1565 ( .A(\gbuff[16][24] ), .B(\gbuff[17][24] ), .C(\gbuff[18][24] ), 
        .D(\gbuff[19][24] ), .S0(n1431), .S1(n1413), .Y(n1313) );
  MX4X1 U1566 ( .A(\gbuff[0][25] ), .B(\gbuff[1][25] ), .C(\gbuff[2][25] ), 
        .D(\gbuff[3][25] ), .S0(n1432), .S1(n1414), .Y(n1327) );
  MX4X1 U1567 ( .A(\gbuff[16][25] ), .B(\gbuff[17][25] ), .C(\gbuff[18][25] ), 
        .D(\gbuff[19][25] ), .S0(n1431), .S1(n1413), .Y(n1323) );
  MX4X1 U1568 ( .A(\gbuff[0][26] ), .B(\gbuff[1][26] ), .C(\gbuff[2][26] ), 
        .D(\gbuff[3][26] ), .S0(n1432), .S1(n1414), .Y(n1337) );
  MX4X1 U1569 ( .A(\gbuff[16][26] ), .B(\gbuff[17][26] ), .C(\gbuff[18][26] ), 
        .D(\gbuff[19][26] ), .S0(n1432), .S1(n1414), .Y(n1333) );
  MX4X1 U1570 ( .A(\gbuff[0][27] ), .B(\gbuff[1][27] ), .C(\gbuff[2][27] ), 
        .D(\gbuff[3][27] ), .S0(n1433), .S1(n1415), .Y(n1347) );
  MX4X1 U1571 ( .A(\gbuff[16][27] ), .B(\gbuff[17][27] ), .C(\gbuff[18][27] ), 
        .D(\gbuff[19][27] ), .S0(n1433), .S1(n1415), .Y(n1343) );
  MX4X1 U1572 ( .A(\gbuff[0][28] ), .B(\gbuff[1][28] ), .C(\gbuff[2][28] ), 
        .D(\gbuff[3][28] ), .S0(n1434), .S1(n1416), .Y(n1357) );
  MX4X1 U1573 ( .A(\gbuff[16][28] ), .B(\gbuff[17][28] ), .C(\gbuff[18][28] ), 
        .D(\gbuff[19][28] ), .S0(n1433), .S1(n1415), .Y(n1353) );
  MX4X1 U1574 ( .A(\gbuff[0][29] ), .B(\gbuff[1][29] ), .C(\gbuff[2][29] ), 
        .D(\gbuff[3][29] ), .S0(n1434), .S1(n1416), .Y(n1367) );
  MX4X1 U1575 ( .A(\gbuff[16][29] ), .B(\gbuff[17][29] ), .C(\gbuff[18][29] ), 
        .D(\gbuff[19][29] ), .S0(n1434), .S1(n1416), .Y(n1363) );
  MX4X1 U1576 ( .A(\gbuff[0][30] ), .B(\gbuff[1][30] ), .C(\gbuff[2][30] ), 
        .D(\gbuff[3][30] ), .S0(n1435), .S1(n1409), .Y(n1377) );
  MX4X1 U1577 ( .A(\gbuff[16][30] ), .B(\gbuff[17][30] ), .C(\gbuff[18][30] ), 
        .D(\gbuff[19][30] ), .S0(n1435), .S1(n1402), .Y(n1373) );
  MX4X1 U1578 ( .A(\gbuff[0][31] ), .B(\gbuff[1][31] ), .C(\gbuff[2][31] ), 
        .D(\gbuff[3][31] ), .S0(n1435), .S1(n1405), .Y(n1387) );
  MX4X1 U1579 ( .A(\gbuff[16][31] ), .B(\gbuff[17][31] ), .C(\gbuff[18][31] ), 
        .D(\gbuff[19][31] ), .S0(n1435), .S1(n1414), .Y(n1383) );
  MX4X1 U1580 ( .A(\gbuff[8][0] ), .B(\gbuff[9][0] ), .C(\gbuff[10][0] ), .D(
        \gbuff[11][0] ), .S0(n1417), .S1(n1398), .Y(n22) );
  MX4X1 U1581 ( .A(\gbuff[24][0] ), .B(\gbuff[25][0] ), .C(\gbuff[26][0] ), 
        .D(\gbuff[27][0] ), .S0(n1437), .S1(n1398), .Y(n18) );
  MX4X1 U1582 ( .A(\gbuff[8][1] ), .B(\gbuff[9][1] ), .C(\gbuff[10][1] ), .D(
        \gbuff[11][1] ), .S0(n1418), .S1(n1399), .Y(n32) );
  MX4X1 U1583 ( .A(\gbuff[24][1] ), .B(\gbuff[25][1] ), .C(\gbuff[26][1] ), 
        .D(\gbuff[27][1] ), .S0(n1418), .S1(n1399), .Y(n28) );
  MX4X1 U1584 ( .A(\gbuff[8][2] ), .B(\gbuff[9][2] ), .C(\gbuff[10][2] ), .D(
        \gbuff[11][2] ), .S0(n1418), .S1(n1399), .Y(n42) );
  MX4X1 U1585 ( .A(\gbuff[24][2] ), .B(\gbuff[25][2] ), .C(\gbuff[26][2] ), 
        .D(\gbuff[27][2] ), .S0(n1418), .S1(n1399), .Y(n38) );
  MX4X1 U1586 ( .A(\gbuff[8][3] ), .B(\gbuff[9][3] ), .C(\gbuff[10][3] ), .D(
        \gbuff[11][3] ), .S0(n1419), .S1(n1400), .Y(n52) );
  MX4X1 U1587 ( .A(\gbuff[24][3] ), .B(\gbuff[25][3] ), .C(\gbuff[26][3] ), 
        .D(\gbuff[27][3] ), .S0(n1419), .S1(n1400), .Y(n48) );
  MX4X1 U1588 ( .A(\gbuff[8][4] ), .B(\gbuff[9][4] ), .C(\gbuff[10][4] ), .D(
        \gbuff[11][4] ), .S0(n1420), .S1(n1401), .Y(n62) );
  MX4X1 U1589 ( .A(\gbuff[24][4] ), .B(\gbuff[25][4] ), .C(\gbuff[26][4] ), 
        .D(\gbuff[27][4] ), .S0(n1419), .S1(n1400), .Y(n58) );
  MX4X1 U1590 ( .A(\gbuff[8][5] ), .B(\gbuff[9][5] ), .C(\gbuff[10][5] ), .D(
        \gbuff[11][5] ), .S0(n1420), .S1(n1401), .Y(n72) );
  MX4X1 U1591 ( .A(\gbuff[24][5] ), .B(\gbuff[25][5] ), .C(\gbuff[26][5] ), 
        .D(\gbuff[27][5] ), .S0(n1420), .S1(n1401), .Y(n68) );
  MX4X1 U1592 ( .A(\gbuff[8][6] ), .B(\gbuff[9][6] ), .C(\gbuff[10][6] ), .D(
        \gbuff[11][6] ), .S0(n1421), .S1(n1402), .Y(n82) );
  MX4X1 U1593 ( .A(\gbuff[24][6] ), .B(\gbuff[25][6] ), .C(\gbuff[26][6] ), 
        .D(\gbuff[27][6] ), .S0(n1421), .S1(n1402), .Y(n78) );
  MX4X1 U1594 ( .A(\gbuff[8][7] ), .B(\gbuff[9][7] ), .C(\gbuff[10][7] ), .D(
        \gbuff[11][7] ), .S0(n1417), .S1(n1403), .Y(n92) );
  MX4X1 U1595 ( .A(\gbuff[24][7] ), .B(\gbuff[25][7] ), .C(\gbuff[26][7] ), 
        .D(\gbuff[27][7] ), .S0(n1421), .S1(n1402), .Y(n88) );
  MX4X1 U1596 ( .A(\gbuff[8][8] ), .B(\gbuff[9][8] ), .C(\gbuff[10][8] ), .D(
        \gbuff[11][8] ), .S0(n1437), .S1(n1403), .Y(n104) );
  MX4X1 U1597 ( .A(\gbuff[24][8] ), .B(\gbuff[25][8] ), .C(\gbuff[26][8] ), 
        .D(\gbuff[27][8] ), .S0(n1436), .S1(n1403), .Y(n98) );
  MX4X1 U1598 ( .A(\gbuff[8][9] ), .B(\gbuff[9][9] ), .C(\gbuff[10][9] ), .D(
        \gbuff[11][9] ), .S0(n1422), .S1(n1404), .Y(n123) );
  MX4X1 U1599 ( .A(\gbuff[24][9] ), .B(\gbuff[25][9] ), .C(\gbuff[26][9] ), 
        .D(\gbuff[27][9] ), .S0(n1436), .S1(n1403), .Y(n116) );
  MX4X1 U1600 ( .A(\gbuff[8][10] ), .B(\gbuff[9][10] ), .C(\gbuff[10][10] ), 
        .D(\gbuff[11][10] ), .S0(n1422), .S1(n1404), .Y(n1175) );
  MX4X1 U1601 ( .A(\gbuff[24][10] ), .B(\gbuff[25][10] ), .C(\gbuff[26][10] ), 
        .D(\gbuff[27][10] ), .S0(n1422), .S1(n1404), .Y(n1171) );
  MX4X1 U1602 ( .A(\gbuff[8][11] ), .B(\gbuff[9][11] ), .C(\gbuff[10][11] ), 
        .D(\gbuff[11][11] ), .S0(n1423), .S1(n1405), .Y(n1185) );
  MX4X1 U1603 ( .A(\gbuff[24][11] ), .B(\gbuff[25][11] ), .C(\gbuff[26][11] ), 
        .D(\gbuff[27][11] ), .S0(n1423), .S1(n1405), .Y(n1181) );
  MX4X1 U1604 ( .A(\gbuff[8][12] ), .B(\gbuff[9][12] ), .C(\gbuff[10][12] ), 
        .D(\gbuff[11][12] ), .S0(n1424), .S1(n1406), .Y(n1195) );
  MX4X1 U1605 ( .A(\gbuff[24][12] ), .B(\gbuff[25][12] ), .C(\gbuff[26][12] ), 
        .D(\gbuff[27][12] ), .S0(n1423), .S1(n1405), .Y(n1191) );
  MX4X1 U1606 ( .A(\gbuff[8][13] ), .B(\gbuff[9][13] ), .C(\gbuff[10][13] ), 
        .D(\gbuff[11][13] ), .S0(n1424), .S1(n1406), .Y(n1205) );
  MX4X1 U1607 ( .A(\gbuff[24][13] ), .B(\gbuff[25][13] ), .C(\gbuff[26][13] ), 
        .D(\gbuff[27][13] ), .S0(n1424), .S1(n1406), .Y(n1201) );
  MX4X1 U1608 ( .A(\gbuff[8][14] ), .B(\gbuff[9][14] ), .C(\gbuff[10][14] ), 
        .D(\gbuff[11][14] ), .S0(n1425), .S1(n1407), .Y(n1215) );
  MX4X1 U1609 ( .A(\gbuff[24][14] ), .B(\gbuff[25][14] ), .C(\gbuff[26][14] ), 
        .D(\gbuff[27][14] ), .S0(n1425), .S1(n1407), .Y(n1211) );
  MX4X1 U1610 ( .A(\gbuff[8][15] ), .B(\gbuff[9][15] ), .C(\gbuff[10][15] ), 
        .D(\gbuff[11][15] ), .S0(n1425), .S1(n1407), .Y(n1225) );
  MX4X1 U1611 ( .A(\gbuff[24][15] ), .B(\gbuff[25][15] ), .C(\gbuff[26][15] ), 
        .D(\gbuff[27][15] ), .S0(n1425), .S1(n1407), .Y(n1221) );
  MX4X1 U1612 ( .A(\gbuff[8][16] ), .B(\gbuff[9][16] ), .C(\gbuff[10][16] ), 
        .D(\gbuff[11][16] ), .S0(n1426), .S1(n1408), .Y(n1235) );
  MX4X1 U1613 ( .A(\gbuff[24][16] ), .B(\gbuff[25][16] ), .C(\gbuff[26][16] ), 
        .D(\gbuff[27][16] ), .S0(n1426), .S1(n1408), .Y(n1231) );
  MX4X1 U1614 ( .A(\gbuff[8][17] ), .B(\gbuff[9][17] ), .C(\gbuff[10][17] ), 
        .D(\gbuff[11][17] ), .S0(n1427), .S1(n1409), .Y(n1245) );
  MX4X1 U1615 ( .A(\gbuff[24][17] ), .B(\gbuff[25][17] ), .C(\gbuff[26][17] ), 
        .D(\gbuff[27][17] ), .S0(n1426), .S1(n1408), .Y(n1241) );
  MX4X1 U1616 ( .A(\gbuff[8][18] ), .B(\gbuff[9][18] ), .C(\gbuff[10][18] ), 
        .D(\gbuff[11][18] ), .S0(n1427), .S1(n1409), .Y(n1255) );
  MX4X1 U1617 ( .A(\gbuff[24][18] ), .B(\gbuff[25][18] ), .C(\gbuff[26][18] ), 
        .D(\gbuff[27][18] ), .S0(n1427), .S1(n1409), .Y(n1251) );
  MX4X1 U1618 ( .A(\gbuff[8][19] ), .B(\gbuff[9][19] ), .C(\gbuff[10][19] ), 
        .D(\gbuff[11][19] ), .S0(n1428), .S1(n1410), .Y(n1265) );
  MX4X1 U1619 ( .A(\gbuff[24][19] ), .B(\gbuff[25][19] ), .C(\gbuff[26][19] ), 
        .D(\gbuff[27][19] ), .S0(n1428), .S1(n1410), .Y(n1261) );
  MX4X1 U1620 ( .A(\gbuff[8][20] ), .B(\gbuff[9][20] ), .C(\gbuff[10][20] ), 
        .D(\gbuff[11][20] ), .S0(n1429), .S1(n1411), .Y(n1275) );
  MX4X1 U1621 ( .A(\gbuff[24][20] ), .B(\gbuff[25][20] ), .C(\gbuff[26][20] ), 
        .D(\gbuff[27][20] ), .S0(n1428), .S1(n1410), .Y(n1271) );
  MX4X1 U1622 ( .A(\gbuff[8][21] ), .B(\gbuff[9][21] ), .C(\gbuff[10][21] ), 
        .D(\gbuff[11][21] ), .S0(n1429), .S1(n1411), .Y(n1285) );
  MX4X1 U1623 ( .A(\gbuff[24][21] ), .B(\gbuff[25][21] ), .C(\gbuff[26][21] ), 
        .D(\gbuff[27][21] ), .S0(n1429), .S1(n1411), .Y(n1281) );
  MX4X1 U1624 ( .A(\gbuff[8][22] ), .B(\gbuff[9][22] ), .C(\gbuff[10][22] ), 
        .D(\gbuff[11][22] ), .S0(n1430), .S1(n1412), .Y(n1295) );
  MX4X1 U1625 ( .A(\gbuff[24][22] ), .B(\gbuff[25][22] ), .C(\gbuff[26][22] ), 
        .D(\gbuff[27][22] ), .S0(n1429), .S1(n1411), .Y(n1291) );
  MX4X1 U1626 ( .A(\gbuff[8][23] ), .B(\gbuff[9][23] ), .C(\gbuff[10][23] ), 
        .D(\gbuff[11][23] ), .S0(n1430), .S1(n1412), .Y(n1305) );
  MX4X1 U1627 ( .A(\gbuff[24][23] ), .B(\gbuff[25][23] ), .C(\gbuff[26][23] ), 
        .D(\gbuff[27][23] ), .S0(n1430), .S1(n1412), .Y(n1301) );
  MX4X1 U1628 ( .A(\gbuff[8][24] ), .B(\gbuff[9][24] ), .C(\gbuff[10][24] ), 
        .D(\gbuff[11][24] ), .S0(n1431), .S1(n1413), .Y(n1315) );
  MX4X1 U1629 ( .A(\gbuff[24][24] ), .B(\gbuff[25][24] ), .C(\gbuff[26][24] ), 
        .D(\gbuff[27][24] ), .S0(n1431), .S1(n1413), .Y(n1311) );
  MX4X1 U1630 ( .A(\gbuff[8][25] ), .B(\gbuff[9][25] ), .C(\gbuff[10][25] ), 
        .D(\gbuff[11][25] ), .S0(n1432), .S1(n1414), .Y(n1325) );
  MX4X1 U1631 ( .A(\gbuff[24][25] ), .B(\gbuff[25][25] ), .C(\gbuff[26][25] ), 
        .D(\gbuff[27][25] ), .S0(n1431), .S1(n1413), .Y(n1321) );
  MX4X1 U1632 ( .A(\gbuff[8][26] ), .B(\gbuff[9][26] ), .C(\gbuff[10][26] ), 
        .D(\gbuff[11][26] ), .S0(n1432), .S1(n1414), .Y(n1335) );
  MX4X1 U1633 ( .A(\gbuff[24][26] ), .B(\gbuff[25][26] ), .C(\gbuff[26][26] ), 
        .D(\gbuff[27][26] ), .S0(n1432), .S1(n1414), .Y(n1331) );
  MX4X1 U1634 ( .A(\gbuff[8][27] ), .B(\gbuff[9][27] ), .C(\gbuff[10][27] ), 
        .D(\gbuff[11][27] ), .S0(n1433), .S1(n1415), .Y(n1345) );
  MX4X1 U1635 ( .A(\gbuff[24][27] ), .B(\gbuff[25][27] ), .C(\gbuff[26][27] ), 
        .D(\gbuff[27][27] ), .S0(n1433), .S1(n1415), .Y(n1341) );
  MX4X1 U1636 ( .A(\gbuff[8][28] ), .B(\gbuff[9][28] ), .C(\gbuff[10][28] ), 
        .D(\gbuff[11][28] ), .S0(n1433), .S1(n1415), .Y(n1355) );
  MX4X1 U1637 ( .A(\gbuff[24][28] ), .B(\gbuff[25][28] ), .C(\gbuff[26][28] ), 
        .D(\gbuff[27][28] ), .S0(n1433), .S1(n1415), .Y(n1351) );
  MX4X1 U1638 ( .A(\gbuff[8][29] ), .B(\gbuff[9][29] ), .C(\gbuff[10][29] ), 
        .D(\gbuff[11][29] ), .S0(n1434), .S1(n1416), .Y(n1365) );
  MX4X1 U1639 ( .A(\gbuff[24][29] ), .B(\gbuff[25][29] ), .C(\gbuff[26][29] ), 
        .D(\gbuff[27][29] ), .S0(n1434), .S1(n1416), .Y(n1361) );
  MX4X1 U1640 ( .A(\gbuff[8][30] ), .B(\gbuff[9][30] ), .C(\gbuff[10][30] ), 
        .D(\gbuff[11][30] ), .S0(n1435), .S1(n1415), .Y(n1375) );
  MX4X1 U1641 ( .A(\gbuff[24][30] ), .B(\gbuff[25][30] ), .C(\gbuff[26][30] ), 
        .D(\gbuff[27][30] ), .S0(n1434), .S1(n1416), .Y(n1371) );
  MX4X1 U1642 ( .A(\gbuff[8][31] ), .B(\gbuff[9][31] ), .C(\gbuff[10][31] ), 
        .D(\gbuff[11][31] ), .S0(n1435), .S1(n1399), .Y(n1385) );
  MX4X1 U1643 ( .A(\gbuff[24][31] ), .B(\gbuff[25][31] ), .C(\gbuff[26][31] ), 
        .D(\gbuff[27][31] ), .S0(n1435), .S1(n1408), .Y(n1381) );
  MX4X1 U1644 ( .A(\gbuff[12][0] ), .B(\gbuff[13][0] ), .C(\gbuff[14][0] ), 
        .D(\gbuff[15][0] ), .S0(n1417), .S1(n1398), .Y(n21) );
  MX4X1 U1645 ( .A(\gbuff[12][1] ), .B(\gbuff[13][1] ), .C(\gbuff[14][1] ), 
        .D(\gbuff[15][1] ), .S0(n1418), .S1(n1399), .Y(n31) );
  MX4X1 U1646 ( .A(\gbuff[12][2] ), .B(\gbuff[13][2] ), .C(\gbuff[14][2] ), 
        .D(\gbuff[15][2] ), .S0(n1418), .S1(n1399), .Y(n41) );
  MX4X1 U1647 ( .A(\gbuff[12][3] ), .B(\gbuff[13][3] ), .C(\gbuff[14][3] ), 
        .D(\gbuff[15][3] ), .S0(n1419), .S1(n1400), .Y(n51) );
  MX4X1 U1648 ( .A(\gbuff[12][4] ), .B(\gbuff[13][4] ), .C(\gbuff[14][4] ), 
        .D(\gbuff[15][4] ), .S0(n1420), .S1(n1401), .Y(n61) );
  MX4X1 U1649 ( .A(\gbuff[12][5] ), .B(\gbuff[13][5] ), .C(\gbuff[14][5] ), 
        .D(\gbuff[15][5] ), .S0(n1420), .S1(n1401), .Y(n71) );
  MX4X1 U1650 ( .A(\gbuff[12][6] ), .B(\gbuff[13][6] ), .C(\gbuff[14][6] ), 
        .D(\gbuff[15][6] ), .S0(n1421), .S1(n1402), .Y(n81) );
  MX4X1 U1651 ( .A(\gbuff[12][7] ), .B(\gbuff[13][7] ), .C(\gbuff[14][7] ), 
        .D(\gbuff[15][7] ), .S0(n1421), .S1(n1402), .Y(n91) );
  MX4X1 U1652 ( .A(\gbuff[12][8] ), .B(\gbuff[13][8] ), .C(\gbuff[14][8] ), 
        .D(\gbuff[15][8] ), .S0(n1437), .S1(n1403), .Y(n101) );
  MX4X1 U1653 ( .A(\gbuff[12][9] ), .B(\gbuff[13][9] ), .C(\gbuff[14][9] ), 
        .D(\gbuff[15][9] ), .S0(n1422), .S1(n1404), .Y(n122) );
  MX4X1 U1654 ( .A(\gbuff[12][10] ), .B(\gbuff[13][10] ), .C(\gbuff[14][10] ), 
        .D(\gbuff[15][10] ), .S0(n1422), .S1(n1404), .Y(n1174) );
  MX4X1 U1655 ( .A(\gbuff[12][11] ), .B(\gbuff[13][11] ), .C(\gbuff[14][11] ), 
        .D(\gbuff[15][11] ), .S0(n1423), .S1(n1405), .Y(n1184) );
  MX4X1 U1656 ( .A(\gbuff[12][12] ), .B(\gbuff[13][12] ), .C(\gbuff[14][12] ), 
        .D(\gbuff[15][12] ), .S0(n1424), .S1(n1406), .Y(n1194) );
  MX4X1 U1657 ( .A(\gbuff[12][13] ), .B(\gbuff[13][13] ), .C(\gbuff[14][13] ), 
        .D(\gbuff[15][13] ), .S0(n1424), .S1(n1406), .Y(n1204) );
  MX4X1 U1658 ( .A(\gbuff[12][14] ), .B(\gbuff[13][14] ), .C(\gbuff[14][14] ), 
        .D(\gbuff[15][14] ), .S0(n1425), .S1(n1407), .Y(n1214) );
  MX4X1 U1659 ( .A(\gbuff[12][15] ), .B(\gbuff[13][15] ), .C(\gbuff[14][15] ), 
        .D(\gbuff[15][15] ), .S0(n1425), .S1(n1407), .Y(n1224) );
  MX4X1 U1660 ( .A(\gbuff[12][16] ), .B(\gbuff[13][16] ), .C(\gbuff[14][16] ), 
        .D(\gbuff[15][16] ), .S0(n1426), .S1(n1408), .Y(n1234) );
  MX4X1 U1661 ( .A(\gbuff[12][17] ), .B(\gbuff[13][17] ), .C(\gbuff[14][17] ), 
        .D(\gbuff[15][17] ), .S0(n1427), .S1(n1409), .Y(n1244) );
  MX4X1 U1662 ( .A(\gbuff[12][18] ), .B(\gbuff[13][18] ), .C(\gbuff[14][18] ), 
        .D(\gbuff[15][18] ), .S0(n1427), .S1(n1409), .Y(n1254) );
  MX4X1 U1663 ( .A(\gbuff[12][19] ), .B(\gbuff[13][19] ), .C(\gbuff[14][19] ), 
        .D(\gbuff[15][19] ), .S0(n1428), .S1(n1410), .Y(n1264) );
  MX4X1 U1664 ( .A(\gbuff[12][20] ), .B(\gbuff[13][20] ), .C(\gbuff[14][20] ), 
        .D(\gbuff[15][20] ), .S0(n1428), .S1(n1410), .Y(n1274) );
  MX4X1 U1665 ( .A(\gbuff[12][21] ), .B(\gbuff[13][21] ), .C(\gbuff[14][21] ), 
        .D(\gbuff[15][21] ), .S0(n1429), .S1(n1411), .Y(n1284) );
  MX4X1 U1666 ( .A(\gbuff[12][22] ), .B(\gbuff[13][22] ), .C(\gbuff[14][22] ), 
        .D(\gbuff[15][22] ), .S0(n1430), .S1(n1412), .Y(n1294) );
  MX4X1 U1667 ( .A(\gbuff[12][23] ), .B(\gbuff[13][23] ), .C(\gbuff[14][23] ), 
        .D(\gbuff[15][23] ), .S0(n1430), .S1(n1412), .Y(n1304) );
  MX4X1 U1668 ( .A(\gbuff[12][24] ), .B(\gbuff[13][24] ), .C(\gbuff[14][24] ), 
        .D(\gbuff[15][24] ), .S0(n1431), .S1(n1413), .Y(n1314) );
  MX4X1 U1669 ( .A(\gbuff[12][25] ), .B(\gbuff[13][25] ), .C(\gbuff[14][25] ), 
        .D(\gbuff[15][25] ), .S0(n1432), .S1(n1414), .Y(n1324) );
  MX4X1 U1670 ( .A(\gbuff[12][26] ), .B(\gbuff[13][26] ), .C(\gbuff[14][26] ), 
        .D(\gbuff[15][26] ), .S0(n1432), .S1(n1414), .Y(n1334) );
  MX4X1 U1671 ( .A(\gbuff[12][27] ), .B(\gbuff[13][27] ), .C(\gbuff[14][27] ), 
        .D(\gbuff[15][27] ), .S0(n1433), .S1(n1415), .Y(n1344) );
  MX4X1 U1672 ( .A(\gbuff[12][28] ), .B(\gbuff[13][28] ), .C(\gbuff[14][28] ), 
        .D(\gbuff[15][28] ), .S0(n1433), .S1(n1415), .Y(n1354) );
  MX4X1 U1673 ( .A(\gbuff[12][29] ), .B(\gbuff[13][29] ), .C(\gbuff[14][29] ), 
        .D(\gbuff[15][29] ), .S0(n1434), .S1(n1416), .Y(n1364) );
  MX4X1 U1674 ( .A(\gbuff[12][30] ), .B(\gbuff[13][30] ), .C(\gbuff[14][30] ), 
        .D(\gbuff[15][30] ), .S0(n1435), .S1(n1398), .Y(n1374) );
  MX4X1 U1675 ( .A(\gbuff[12][31] ), .B(\gbuff[13][31] ), .C(\gbuff[14][31] ), 
        .D(\gbuff[15][31] ), .S0(n1435), .S1(n1398), .Y(n1384) );
  MXI2X1 U1676 ( .A(n25), .B(n26), .S0(n1390), .Y(N47) );
  MXI4X1 U1677 ( .A(n20), .B(n18), .C(n19), .D(n17), .S0(n1393), .S1(n1395), 
        .Y(n26) );
  MXI4X1 U1678 ( .A(n24), .B(n22), .C(n23), .D(n21), .S0(n1394), .S1(n1395), 
        .Y(n25) );
  MX4X1 U1679 ( .A(\gbuff[28][0] ), .B(\gbuff[29][0] ), .C(\gbuff[30][0] ), 
        .D(\gbuff[31][0] ), .S0(n1437), .S1(n1398), .Y(n17) );
  MXI2X1 U1680 ( .A(n35), .B(n36), .S0(n1390), .Y(N46) );
  MXI4X1 U1681 ( .A(n30), .B(n28), .C(n29), .D(n27), .S0(n1394), .S1(n1396), 
        .Y(n36) );
  MXI4X1 U1682 ( .A(n34), .B(n32), .C(n33), .D(n31), .S0(n1392), .S1(n1397), 
        .Y(n35) );
  MX4X1 U1683 ( .A(\gbuff[28][1] ), .B(\gbuff[29][1] ), .C(\gbuff[30][1] ), 
        .D(\gbuff[31][1] ), .S0(n1437), .S1(n1398), .Y(n27) );
  MXI2X1 U1684 ( .A(n45), .B(n46), .S0(n1390), .Y(N45) );
  MXI4X1 U1685 ( .A(n40), .B(n38), .C(n39), .D(n37), .S0(n1391), .S1(n1395), 
        .Y(n46) );
  MXI4X1 U1686 ( .A(n44), .B(n42), .C(n43), .D(n41), .S0(n1391), .S1(n1395), 
        .Y(n45) );
  MX4X1 U1687 ( .A(\gbuff[28][2] ), .B(\gbuff[29][2] ), .C(\gbuff[30][2] ), 
        .D(\gbuff[31][2] ), .S0(n1418), .S1(n1399), .Y(n37) );
  MXI2X1 U1688 ( .A(n55), .B(n56), .S0(n1390), .Y(N44) );
  MXI4X1 U1689 ( .A(n50), .B(n48), .C(n49), .D(n47), .S0(n1391), .S1(n1395), 
        .Y(n56) );
  MXI4X1 U1690 ( .A(n54), .B(n52), .C(n53), .D(n51), .S0(n1391), .S1(n1395), 
        .Y(n55) );
  MX4X1 U1691 ( .A(\gbuff[28][3] ), .B(\gbuff[29][3] ), .C(\gbuff[30][3] ), 
        .D(\gbuff[31][3] ), .S0(n1419), .S1(n1400), .Y(n47) );
  MXI2X1 U1692 ( .A(n65), .B(n66), .S0(n1390), .Y(N43) );
  MXI4X1 U1693 ( .A(n60), .B(n58), .C(n59), .D(n57), .S0(n1391), .S1(n1395), 
        .Y(n66) );
  MXI4X1 U1694 ( .A(n64), .B(n62), .C(n63), .D(n61), .S0(n1391), .S1(n1395), 
        .Y(n65) );
  MX4X1 U1695 ( .A(\gbuff[28][4] ), .B(\gbuff[29][4] ), .C(\gbuff[30][4] ), 
        .D(\gbuff[31][4] ), .S0(n1419), .S1(n1400), .Y(n57) );
  MXI2X1 U1696 ( .A(n75), .B(n76), .S0(n1738), .Y(N42) );
  MXI4X1 U1697 ( .A(n70), .B(n68), .C(n69), .D(n67), .S0(n1391), .S1(n1395), 
        .Y(n76) );
  MXI4X1 U1698 ( .A(n74), .B(n72), .C(n73), .D(n71), .S0(n1391), .S1(n1395), 
        .Y(n75) );
  MX4X1 U1699 ( .A(\gbuff[28][5] ), .B(\gbuff[29][5] ), .C(\gbuff[30][5] ), 
        .D(\gbuff[31][5] ), .S0(n1420), .S1(n1401), .Y(n67) );
  MXI2X1 U1700 ( .A(n85), .B(n86), .S0(n1390), .Y(N41) );
  MXI4X1 U1701 ( .A(n80), .B(n78), .C(n79), .D(n77), .S0(n1391), .S1(n1395), 
        .Y(n86) );
  MXI4X1 U1702 ( .A(n84), .B(n82), .C(n83), .D(n81), .S0(n1391), .S1(n1395), 
        .Y(n85) );
  MX4X1 U1703 ( .A(\gbuff[28][6] ), .B(\gbuff[29][6] ), .C(\gbuff[30][6] ), 
        .D(\gbuff[31][6] ), .S0(n1421), .S1(n1402), .Y(n77) );
  MXI2X1 U1704 ( .A(n95), .B(n96), .S0(n1738), .Y(N40) );
  MXI4X1 U1705 ( .A(n90), .B(n88), .C(n89), .D(n87), .S0(n1391), .S1(n1395), 
        .Y(n96) );
  MXI4X1 U1706 ( .A(n94), .B(n92), .C(n93), .D(n91), .S0(n1391), .S1(n1395), 
        .Y(n95) );
  MX4X1 U1707 ( .A(\gbuff[28][7] ), .B(\gbuff[29][7] ), .C(\gbuff[30][7] ), 
        .D(\gbuff[31][7] ), .S0(n1421), .S1(n1402), .Y(n87) );
  MXI2X1 U1708 ( .A(n110), .B(n112), .S0(n1390), .Y(N39) );
  MXI4X1 U1709 ( .A(n100), .B(n98), .C(n99), .D(n97), .S0(n1393), .S1(n1396), 
        .Y(n112) );
  MXI4X1 U1710 ( .A(n108), .B(n104), .C(n106), .D(n101), .S0(n1392), .S1(n1396), .Y(n110) );
  MX4X1 U1711 ( .A(\gbuff[28][8] ), .B(\gbuff[29][8] ), .C(\gbuff[30][8] ), 
        .D(\gbuff[31][8] ), .S0(n1436), .S1(n1403), .Y(n97) );
  MXI2X1 U1712 ( .A(n126), .B(n127), .S0(n1390), .Y(N38) );
  MXI4X1 U1713 ( .A(n121), .B(n116), .C(n119), .D(n114), .S0(n1394), .S1(n1396), .Y(n127) );
  MXI4X1 U1714 ( .A(n125), .B(n123), .C(n124), .D(n122), .S0(n1393), .S1(n1396), .Y(n126) );
  MX4X1 U1715 ( .A(\gbuff[28][9] ), .B(\gbuff[29][9] ), .C(\gbuff[30][9] ), 
        .D(\gbuff[31][9] ), .S0(n1437), .S1(n1403), .Y(n114) );
  MXI2X1 U1716 ( .A(n1178), .B(n1179), .S0(n1390), .Y(N37) );
  MXI4X1 U1717 ( .A(n1173), .B(n1171), .C(n1172), .D(n1170), .S0(n1391), .S1(
        n1396), .Y(n1179) );
  MXI4X1 U1718 ( .A(n1177), .B(n1175), .C(n1176), .D(n1174), .S0(n1392), .S1(
        n1396), .Y(n1178) );
  MX4X1 U1719 ( .A(\gbuff[28][10] ), .B(\gbuff[29][10] ), .C(\gbuff[30][10] ), 
        .D(\gbuff[31][10] ), .S0(n1422), .S1(n1404), .Y(n1170) );
  MXI2X1 U1720 ( .A(n1188), .B(n1189), .S0(n1390), .Y(N36) );
  MXI4X1 U1721 ( .A(n1183), .B(n1181), .C(n1182), .D(n1180), .S0(n1391), .S1(
        n1396), .Y(n1189) );
  MXI4X1 U1722 ( .A(n1187), .B(n1185), .C(n1186), .D(n1184), .S0(n1393), .S1(
        n1396), .Y(n1188) );
  MX4X1 U1723 ( .A(\gbuff[28][11] ), .B(\gbuff[29][11] ), .C(\gbuff[30][11] ), 
        .D(\gbuff[31][11] ), .S0(n1423), .S1(n1405), .Y(n1180) );
  MXI2X1 U1724 ( .A(n1198), .B(n1199), .S0(n1390), .Y(N35) );
  MXI4X1 U1725 ( .A(n1193), .B(n1191), .C(n1192), .D(n1190), .S0(n1391), .S1(
        n1396), .Y(n1199) );
  MXI4X1 U1726 ( .A(n1197), .B(n1195), .C(n1196), .D(n1194), .S0(n1394), .S1(
        n1396), .Y(n1198) );
  MX4X1 U1727 ( .A(\gbuff[28][12] ), .B(\gbuff[29][12] ), .C(\gbuff[30][12] ), 
        .D(\gbuff[31][12] ), .S0(n1423), .S1(n1405), .Y(n1190) );
  MXI2X1 U1728 ( .A(n1208), .B(n1209), .S0(n1390), .Y(N34) );
  MXI4X1 U1729 ( .A(n1203), .B(n1201), .C(n1202), .D(n1200), .S0(n1391), .S1(
        n1396), .Y(n1209) );
  MXI4X1 U1730 ( .A(n1207), .B(n1205), .C(n1206), .D(n1204), .S0(n1392), .S1(
        n1396), .Y(n1208) );
  MX4X1 U1731 ( .A(\gbuff[28][13] ), .B(\gbuff[29][13] ), .C(\gbuff[30][13] ), 
        .D(\gbuff[31][13] ), .S0(n1424), .S1(n1406), .Y(n1200) );
  MXI2X1 U1732 ( .A(n1218), .B(n1219), .S0(n1390), .Y(N33) );
  MXI4X1 U1733 ( .A(n1213), .B(n1211), .C(n1212), .D(n1210), .S0(n1392), .S1(
        n1397), .Y(n1219) );
  MXI4X1 U1734 ( .A(n1217), .B(n1215), .C(n1216), .D(n1214), .S0(n1392), .S1(
        n1396), .Y(n1218) );
  MX4X1 U1735 ( .A(\gbuff[28][14] ), .B(\gbuff[29][14] ), .C(\gbuff[30][14] ), 
        .D(\gbuff[31][14] ), .S0(n1424), .S1(n1406), .Y(n1210) );
  MXI2X1 U1736 ( .A(n1228), .B(n1229), .S0(n1390), .Y(N32) );
  MXI4X1 U1737 ( .A(n1223), .B(n1221), .C(n1222), .D(n1220), .S0(n1392), .S1(
        n1396), .Y(n1229) );
  MXI4X1 U1738 ( .A(n1227), .B(n1225), .C(n1226), .D(n1224), .S0(n1392), .S1(
        n1396), .Y(n1228) );
  MX4X1 U1739 ( .A(\gbuff[28][15] ), .B(\gbuff[29][15] ), .C(\gbuff[30][15] ), 
        .D(\gbuff[31][15] ), .S0(n1425), .S1(n1407), .Y(n1220) );
  MXI2X1 U1740 ( .A(n1238), .B(n1239), .S0(n1390), .Y(N31) );
  MXI4X1 U1741 ( .A(n1233), .B(n1231), .C(n1232), .D(n1230), .S0(n1392), .S1(
        n1395), .Y(n1239) );
  MXI4X1 U1742 ( .A(n1237), .B(n1235), .C(n1236), .D(n1234), .S0(n1392), .S1(
        n1397), .Y(n1238) );
  MX4X1 U1743 ( .A(\gbuff[28][16] ), .B(\gbuff[29][16] ), .C(\gbuff[30][16] ), 
        .D(\gbuff[31][16] ), .S0(n1426), .S1(n1408), .Y(n1230) );
  MXI2X1 U1744 ( .A(n1248), .B(n1249), .S0(n1390), .Y(N30) );
  MXI4X1 U1745 ( .A(n1243), .B(n1241), .C(n1242), .D(n1240), .S0(n1392), .S1(
        n1396), .Y(n1249) );
  MXI4X1 U1746 ( .A(n1247), .B(n1245), .C(n1246), .D(n1244), .S0(n1392), .S1(
        n1396), .Y(n1248) );
  MX4X1 U1747 ( .A(\gbuff[28][17] ), .B(\gbuff[29][17] ), .C(\gbuff[30][17] ), 
        .D(\gbuff[31][17] ), .S0(n1426), .S1(n1408), .Y(n1240) );
  MXI2X1 U1748 ( .A(n1258), .B(n1259), .S0(n1390), .Y(N29) );
  MXI4X1 U1749 ( .A(n1253), .B(n1251), .C(n1252), .D(n1250), .S0(n1392), .S1(
        n1397), .Y(n1259) );
  MXI4X1 U1750 ( .A(n1257), .B(n1255), .C(n1256), .D(n1254), .S0(n1392), .S1(
        n1395), .Y(n1258) );
  MX4X1 U1751 ( .A(\gbuff[28][18] ), .B(\gbuff[29][18] ), .C(\gbuff[30][18] ), 
        .D(\gbuff[31][18] ), .S0(n1427), .S1(n1409), .Y(n1250) );
  MXI2X1 U1752 ( .A(n1268), .B(n1269), .S0(n1390), .Y(N28) );
  MXI4X1 U1753 ( .A(n1263), .B(n1261), .C(n1262), .D(n1260), .S0(n1392), .S1(
        n1396), .Y(n1269) );
  MXI4X1 U1754 ( .A(n1267), .B(n1265), .C(n1266), .D(n1264), .S0(n1392), .S1(
        n1396), .Y(n1268) );
  MX4X1 U1755 ( .A(\gbuff[28][19] ), .B(\gbuff[29][19] ), .C(\gbuff[30][19] ), 
        .D(\gbuff[31][19] ), .S0(n1428), .S1(n1410), .Y(n1260) );
  MXI2X1 U1756 ( .A(n1278), .B(n1279), .S0(n1738), .Y(N27) );
  MXI4X1 U1757 ( .A(n1273), .B(n1271), .C(n1272), .D(n1270), .S0(n1393), .S1(
        n1397), .Y(n1279) );
  MXI4X1 U1758 ( .A(n1277), .B(n1275), .C(n1276), .D(n1274), .S0(n1393), .S1(
        n1397), .Y(n1278) );
  MX4X1 U1759 ( .A(\gbuff[28][20] ), .B(\gbuff[29][20] ), .C(\gbuff[30][20] ), 
        .D(\gbuff[31][20] ), .S0(n1428), .S1(n1410), .Y(n1270) );
  MXI2X1 U1760 ( .A(n1288), .B(n1289), .S0(N14), .Y(N26) );
  MXI4X1 U1761 ( .A(n1283), .B(n1281), .C(n1282), .D(n1280), .S0(n1393), .S1(
        n1397), .Y(n1289) );
  MXI4X1 U1762 ( .A(n1287), .B(n1285), .C(n1286), .D(n1284), .S0(n1393), .S1(
        n1397), .Y(n1288) );
  MX4X1 U1763 ( .A(\gbuff[28][21] ), .B(\gbuff[29][21] ), .C(\gbuff[30][21] ), 
        .D(\gbuff[31][21] ), .S0(n1429), .S1(n1411), .Y(n1280) );
  MXI2X1 U1764 ( .A(n1298), .B(n1299), .S0(N14), .Y(N25) );
  MXI4X1 U1765 ( .A(n1293), .B(n1291), .C(n1292), .D(n1290), .S0(n1393), .S1(
        n1397), .Y(n1299) );
  MXI4X1 U1766 ( .A(n1297), .B(n1295), .C(n1296), .D(n1294), .S0(n1393), .S1(
        n1397), .Y(n1298) );
  MX4X1 U1767 ( .A(\gbuff[28][22] ), .B(\gbuff[29][22] ), .C(\gbuff[30][22] ), 
        .D(\gbuff[31][22] ), .S0(n1429), .S1(n1411), .Y(n1290) );
  MXI2X1 U1768 ( .A(n1308), .B(n1309), .S0(N14), .Y(N24) );
  MXI4X1 U1769 ( .A(n1303), .B(n1301), .C(n1302), .D(n1300), .S0(n1393), .S1(
        n1397), .Y(n1309) );
  MXI4X1 U1770 ( .A(n1307), .B(n1305), .C(n1306), .D(n1304), .S0(n1393), .S1(
        n1397), .Y(n1308) );
  MX4X1 U1771 ( .A(\gbuff[28][23] ), .B(\gbuff[29][23] ), .C(\gbuff[30][23] ), 
        .D(\gbuff[31][23] ), .S0(n1430), .S1(n1412), .Y(n1300) );
  MXI2X1 U1772 ( .A(n1318), .B(n1319), .S0(N14), .Y(N23) );
  MXI4X1 U1773 ( .A(n1313), .B(n1311), .C(n1312), .D(n1310), .S0(n1393), .S1(
        n1397), .Y(n1319) );
  MXI4X1 U1774 ( .A(n1317), .B(n1315), .C(n1316), .D(n1314), .S0(n1393), .S1(
        n1397), .Y(n1318) );
  MX4X1 U1775 ( .A(\gbuff[28][24] ), .B(\gbuff[29][24] ), .C(\gbuff[30][24] ), 
        .D(\gbuff[31][24] ), .S0(n1431), .S1(n1413), .Y(n1310) );
  MXI2X1 U1776 ( .A(n1328), .B(n1329), .S0(N14), .Y(N22) );
  MXI4X1 U1777 ( .A(n1323), .B(n1321), .C(n1322), .D(n1320), .S0(n1393), .S1(
        n1397), .Y(n1329) );
  MXI4X1 U1778 ( .A(n1327), .B(n1325), .C(n1326), .D(n1324), .S0(n1393), .S1(
        n1397), .Y(n1328) );
  MX4X1 U1779 ( .A(\gbuff[28][25] ), .B(\gbuff[29][25] ), .C(\gbuff[30][25] ), 
        .D(\gbuff[31][25] ), .S0(n1431), .S1(n1413), .Y(n1320) );
  MXI2X1 U1780 ( .A(n1338), .B(n1339), .S0(n1738), .Y(N21) );
  MXI4X1 U1781 ( .A(n1333), .B(n1331), .C(n1332), .D(n1330), .S0(n1394), .S1(
        n1397), .Y(n1339) );
  MXI4X1 U1782 ( .A(n1337), .B(n1335), .C(n1336), .D(n1334), .S0(n1394), .S1(
        n1397), .Y(n1338) );
  MX4X1 U1783 ( .A(\gbuff[28][26] ), .B(\gbuff[29][26] ), .C(\gbuff[30][26] ), 
        .D(\gbuff[31][26] ), .S0(n1432), .S1(n1414), .Y(n1330) );
  MXI2X1 U1784 ( .A(n1348), .B(n1349), .S0(n1738), .Y(N20) );
  MXI4X1 U1785 ( .A(n1343), .B(n1341), .C(n1342), .D(n1340), .S0(n1394), .S1(
        n1395), .Y(n1349) );
  MXI4X1 U1786 ( .A(n1347), .B(n1345), .C(n1346), .D(n1344), .S0(n1394), .S1(
        n1395), .Y(n1348) );
  MX4X1 U1787 ( .A(\gbuff[28][27] ), .B(\gbuff[29][27] ), .C(\gbuff[30][27] ), 
        .D(\gbuff[31][27] ), .S0(n1432), .S1(n1414), .Y(n1340) );
  MXI2X1 U1788 ( .A(n1358), .B(n1359), .S0(n1738), .Y(N19) );
  MXI4X1 U1789 ( .A(n1353), .B(n1351), .C(n1352), .D(n1350), .S0(n1394), .S1(
        n1735), .Y(n1359) );
  MXI4X1 U1790 ( .A(n1357), .B(n1355), .C(n1356), .D(n1354), .S0(n1394), .S1(
        n1397), .Y(n1358) );
  MX4X1 U1791 ( .A(\gbuff[28][28] ), .B(\gbuff[29][28] ), .C(\gbuff[30][28] ), 
        .D(\gbuff[31][28] ), .S0(n1433), .S1(n1415), .Y(n1350) );
  MXI2X1 U1792 ( .A(n1368), .B(n1369), .S0(n1738), .Y(N18) );
  MXI4X1 U1793 ( .A(n1363), .B(n1361), .C(n1362), .D(n1360), .S0(n1394), .S1(
        N12), .Y(n1369) );
  MXI4X1 U1794 ( .A(n1367), .B(n1365), .C(n1366), .D(n1364), .S0(n1394), .S1(
        n1395), .Y(n1368) );
  MX4X1 U1795 ( .A(\gbuff[28][29] ), .B(\gbuff[29][29] ), .C(\gbuff[30][29] ), 
        .D(\gbuff[31][29] ), .S0(n1434), .S1(n1416), .Y(n1360) );
  MXI2X1 U1796 ( .A(n1378), .B(n1379), .S0(n1738), .Y(N17) );
  MXI4X1 U1797 ( .A(n1373), .B(n1371), .C(n1372), .D(n1370), .S0(n1394), .S1(
        N12), .Y(n1379) );
  MXI4X1 U1798 ( .A(n1377), .B(n1375), .C(n1376), .D(n1374), .S0(n1394), .S1(
        n1397), .Y(n1378) );
  MX4X1 U1799 ( .A(\gbuff[28][30] ), .B(\gbuff[29][30] ), .C(\gbuff[30][30] ), 
        .D(\gbuff[31][30] ), .S0(n1434), .S1(n1416), .Y(n1370) );
  MXI2X1 U1800 ( .A(n1388), .B(n1389), .S0(n1738), .Y(N16) );
  MXI4X1 U1801 ( .A(n1383), .B(n1381), .C(n1382), .D(n1380), .S0(n1394), .S1(
        N12), .Y(n1389) );
  MXI4X1 U1802 ( .A(n1387), .B(n1385), .C(n1386), .D(n1384), .S0(n1394), .S1(
        n1395), .Y(n1388) );
  MX4X1 U1803 ( .A(\gbuff[28][31] ), .B(\gbuff[29][31] ), .C(\gbuff[30][31] ), 
        .D(\gbuff[31][31] ), .S0(n1435), .S1(n1416), .Y(n1380) );
  CLKBUFX3 U1804 ( .A(N12), .Y(n1735) );
  CLKBUFX3 U1805 ( .A(N14), .Y(n1738) );
endmodule


module pe_0_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U85 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U86 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U87 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U91 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(a[5]), .Y(n123) );
  CLKINVX1 U95 ( .A(b[5]), .Y(n129) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_0 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_0_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, N3, N2, N1}) );
  pe_0_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_15_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U85 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U86 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U87 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U91 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(a[5]), .Y(n123) );
  CLKINVX1 U95 ( .A(b[5]), .Y(n129) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_15_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_15 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_15_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, 
        N3, N2, N1}) );
  pe_15_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_14_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U85 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U86 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U87 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U91 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(a[5]), .Y(n123) );
  CLKINVX1 U95 ( .A(b[5]), .Y(n129) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_14_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_14 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_14_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, 
        N3, N2, N1}) );
  pe_14_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_13_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U85 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U86 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U87 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U91 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(a[5]), .Y(n123) );
  CLKINVX1 U95 ( .A(b[5]), .Y(n129) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_13_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_13 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_13_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, 
        N3, N2, N1}) );
  pe_13_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_12_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U85 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U86 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U87 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U91 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(a[5]), .Y(n123) );
  CLKINVX1 U95 ( .A(b[5]), .Y(n129) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_12_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_12 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_12_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, 
        N3, N2, N1}) );
  pe_12_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_11_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U85 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U86 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U87 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U91 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(a[5]), .Y(n123) );
  CLKINVX1 U95 ( .A(b[5]), .Y(n129) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_11_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_11 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_11_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, 
        N3, N2, N1}) );
  pe_11_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_10_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U85 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U86 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U87 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U91 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(b[5]), .Y(n129) );
  CLKINVX1 U95 ( .A(a[5]), .Y(n123) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_10_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_10 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_10_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, 
        N3, N2, N1}) );
  pe_10_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_9_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U85 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U86 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U87 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U91 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(b[5]), .Y(n129) );
  CLKINVX1 U95 ( .A(a[5]), .Y(n123) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_9_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_9 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_9_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, N3, N2, N1}) );
  pe_9_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_8_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U85 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U86 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U87 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U91 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(a[5]), .Y(n123) );
  CLKINVX1 U95 ( .A(b[5]), .Y(n129) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_8_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_8 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_8_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, N3, N2, N1}) );
  pe_8_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_7_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U85 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U86 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U87 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U91 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(b[5]), .Y(n129) );
  CLKINVX1 U95 ( .A(a[5]), .Y(n123) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_7_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_7 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_7_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, N3, N2, N1}) );
  pe_7_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_6_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U85 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U86 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U87 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U91 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(b[5]), .Y(n129) );
  CLKINVX1 U95 ( .A(a[5]), .Y(n123) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_6_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_6 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_6_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, N3, N2, N1}) );
  pe_6_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_5_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U85 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U86 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U87 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U91 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(a[5]), .Y(n123) );
  CLKINVX1 U95 ( .A(b[5]), .Y(n129) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_5_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_5 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_5_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, N3, N2, N1}) );
  pe_5_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_4_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U85 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U86 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U87 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U91 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(a[5]), .Y(n123) );
  CLKINVX1 U95 ( .A(b[5]), .Y(n129) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_4_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_4 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_4_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, N3, N2, N1}) );
  pe_4_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_3_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U85 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U86 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U87 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U91 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(b[5]), .Y(n129) );
  CLKINVX1 U95 ( .A(a[5]), .Y(n123) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_3_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_3 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_3_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, N3, N2, N1}) );
  pe_3_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_2_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U85 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U86 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U87 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U91 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(a[5]), .Y(n123) );
  CLKINVX1 U95 ( .A(b[5]), .Y(n129) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_2 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_2_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, N3, N2, N1}) );
  pe_2_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module pe_1_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n46, n48, n49, n51, n52, n53, n55, n56, n57, n58, n60,
         n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  ADDFXL U3 ( .A(n20), .B(n27), .CI(n3), .CO(n2), .S(product[6]) );
  ADDFXL U4 ( .A(n28), .B(n34), .CI(n4), .CO(n3), .S(product[5]) );
  ADDFXL U5 ( .A(n35), .B(n38), .CI(n5), .CO(n4), .S(product[4]) );
  ADDFXL U6 ( .A(n39), .B(n41), .CI(n6), .CO(n5), .S(product[3]) );
  ADDFXL U7 ( .A(n7), .B(n64), .CI(n43), .CO(n6), .S(product[2]) );
  ADDHXL U8 ( .A(n71), .B(n78), .CO(n7), .S(product[1]) );
  CMPR42X1 U19 ( .A(n60), .B(n25), .C(n26), .D(n29), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  CMPR42X1 U20 ( .A(n73), .B(n51), .C(n66), .D(n55), .ICI(n31), .S(n23), .ICO(
        n21), .CO(n22) );
  ADDHXL U21 ( .A(n48), .B(n46), .CO(n24), .S(n25) );
  CMPR42X1 U22 ( .A(n67), .B(n36), .C(n33), .D(n32), .ICI(n30), .S(n28), .ICO(
        n26), .CO(n27) );
  ADDFXL U23 ( .A(n56), .B(n74), .CI(n61), .CO(n29), .S(n30) );
  ADDHXL U24 ( .A(n52), .B(n49), .CO(n31), .S(n32) );
  CMPR42X1 U25 ( .A(n75), .B(n62), .C(n68), .D(n40), .ICI(n37), .S(n35), .ICO(
        n33), .CO(n34) );
  ADDHXL U26 ( .A(n57), .B(n53), .CO(n36), .S(n37) );
  ADDFXL U27 ( .A(n69), .B(n76), .CI(n42), .CO(n38), .S(n39) );
  ADDHXL U28 ( .A(n63), .B(n58), .CO(n40), .S(n41) );
  ADDHXL U29 ( .A(n77), .B(n70), .CO(n42), .S(n43) );
  CLKINVX1 U84 ( .A(a[1]), .Y(n127) );
  CLKINVX1 U85 ( .A(b[0]), .Y(n134) );
  CLKINVX1 U86 ( .A(a[0]), .Y(n128) );
  CLKINVX1 U87 ( .A(b[1]), .Y(n133) );
  CLKINVX1 U88 ( .A(b[2]), .Y(n132) );
  CLKINVX1 U89 ( .A(a[2]), .Y(n126) );
  CLKINVX1 U90 ( .A(a[3]), .Y(n125) );
  CLKINVX1 U91 ( .A(b[3]), .Y(n131) );
  CLKINVX1 U92 ( .A(a[4]), .Y(n124) );
  CLKINVX1 U93 ( .A(b[4]), .Y(n130) );
  CLKINVX1 U94 ( .A(a[5]), .Y(n123) );
  CLKINVX1 U95 ( .A(b[5]), .Y(n129) );
  XOR2X1 U96 ( .A(n135), .B(n136), .Y(product[7]) );
  XOR2X1 U97 ( .A(n137), .B(n138), .Y(n136) );
  XOR2X1 U98 ( .A(n139), .B(n140), .Y(n138) );
  NAND2X1 U99 ( .A(b[5]), .B(a[2]), .Y(n140) );
  NAND2X1 U100 ( .A(b[4]), .B(a[3]), .Y(n139) );
  XOR2X1 U101 ( .A(n141), .B(n142), .Y(n137) );
  XOR2X1 U102 ( .A(n143), .B(n144), .Y(n142) );
  XOR2X1 U103 ( .A(n145), .B(n146), .Y(n144) );
  NAND2X1 U104 ( .A(b[3]), .B(a[4]), .Y(n146) );
  NAND2X1 U105 ( .A(b[2]), .B(a[5]), .Y(n145) );
  XOR2X1 U106 ( .A(n147), .B(n148), .Y(n143) );
  NAND2X1 U107 ( .A(b[7]), .B(a[0]), .Y(n148) );
  NAND2X1 U108 ( .A(b[1]), .B(a[6]), .Y(n147) );
  XOR2X1 U109 ( .A(n149), .B(n150), .Y(n141) );
  XOR2X1 U110 ( .A(n151), .B(n18), .Y(n150) );
  NAND2X1 U111 ( .A(b[0]), .B(a[7]), .Y(n151) );
  XNOR2X1 U112 ( .A(n22), .B(n19), .Y(n149) );
  XOR2X1 U113 ( .A(n152), .B(n153), .Y(n135) );
  XOR2X1 U114 ( .A(n154), .B(n2), .Y(n153) );
  NAND2X1 U115 ( .A(b[6]), .B(a[1]), .Y(n154) );
  XNOR2X1 U116 ( .A(n24), .B(n21), .Y(n152) );
  NOR2X1 U117 ( .A(n134), .B(n128), .Y(product[0]) );
  NOR2X1 U118 ( .A(n133), .B(n128), .Y(n78) );
  NOR2X1 U119 ( .A(n128), .B(n132), .Y(n77) );
  NOR2X1 U120 ( .A(n128), .B(n131), .Y(n76) );
  NOR2X1 U121 ( .A(n128), .B(n130), .Y(n75) );
  NOR2X1 U122 ( .A(n128), .B(n129), .Y(n74) );
  AND2X1 U123 ( .A(b[6]), .B(a[0]), .Y(n73) );
  NOR2X1 U124 ( .A(n127), .B(n134), .Y(n71) );
  NOR2X1 U125 ( .A(n127), .B(n133), .Y(n70) );
  NOR2X1 U126 ( .A(n127), .B(n132), .Y(n69) );
  NOR2X1 U127 ( .A(n127), .B(n131), .Y(n68) );
  NOR2X1 U128 ( .A(n127), .B(n130), .Y(n67) );
  NOR2X1 U129 ( .A(n127), .B(n129), .Y(n66) );
  NOR2X1 U130 ( .A(n134), .B(n126), .Y(n64) );
  NOR2X1 U131 ( .A(n133), .B(n126), .Y(n63) );
  NOR2X1 U132 ( .A(n132), .B(n126), .Y(n62) );
  NOR2X1 U133 ( .A(n131), .B(n126), .Y(n61) );
  NOR2X1 U134 ( .A(n130), .B(n126), .Y(n60) );
  NOR2X1 U135 ( .A(n134), .B(n125), .Y(n58) );
  NOR2X1 U136 ( .A(n133), .B(n125), .Y(n57) );
  NOR2X1 U137 ( .A(n132), .B(n125), .Y(n56) );
  NOR2X1 U138 ( .A(n131), .B(n125), .Y(n55) );
  NOR2X1 U139 ( .A(n134), .B(n124), .Y(n53) );
  NOR2X1 U140 ( .A(n133), .B(n124), .Y(n52) );
  NOR2X1 U141 ( .A(n132), .B(n124), .Y(n51) );
  NOR2X1 U142 ( .A(n134), .B(n123), .Y(n49) );
  NOR2X1 U143 ( .A(n133), .B(n123), .Y(n48) );
  AND2X1 U144 ( .A(a[6]), .B(b[0]), .Y(n46) );
endmodule


module pe_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module pe_1 ( clk, rst, a, b, psum, a_out, out );
  input [7:0] a;
  input [7:0] b;
  input [7:0] psum;
  output [7:0] a_out;
  output [7:0] out;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N8, N7, N6, N5, N4, N3, N2, N1,
         n1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  pe_1_DW_mult_uns_0 mult_19 ( .a(a), .b(b), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, N8, N7, N6, N5, N4, N3, N2, N1}) );
  pe_1_DW01_add_0 add_19 ( .A({N8, N7, N6, N5, N4, N3, N2, N1}), .B(psum), 
        .CI(1'b0), .SUM({N16, N15, N14, N13, N12, N11, N10, N9}) );
  DFFRX1 \out_reg[7]  ( .D(N16), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFRX1 \out_reg[6]  ( .D(N15), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFRX1 \out_reg[5]  ( .D(N14), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFRX1 \out_reg[4]  ( .D(N13), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFRX1 \out_reg[3]  ( .D(N12), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFRX1 \out_reg[2]  ( .D(N11), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFRX1 \out_reg[1]  ( .D(N10), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFRX1 \out_reg[0]  ( .D(N9), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFRX1 \a_out_reg[7]  ( .D(a[7]), .CK(clk), .RN(n1), .Q(a_out[7]) );
  DFFRX1 \a_out_reg[6]  ( .D(a[6]), .CK(clk), .RN(n1), .Q(a_out[6]) );
  DFFRX1 \a_out_reg[5]  ( .D(a[5]), .CK(clk), .RN(n1), .Q(a_out[5]) );
  DFFRX1 \a_out_reg[4]  ( .D(a[4]), .CK(clk), .RN(n1), .Q(a_out[4]) );
  DFFRX1 \a_out_reg[3]  ( .D(a[3]), .CK(clk), .RN(n1), .Q(a_out[3]) );
  DFFRX1 \a_out_reg[2]  ( .D(a[2]), .CK(clk), .RN(n1), .Q(a_out[2]) );
  DFFRX1 \a_out_reg[1]  ( .D(a[1]), .CK(clk), .RN(n1), .Q(a_out[1]) );
  DFFRX1 \a_out_reg[0]  ( .D(a[0]), .CK(clk), .RN(n1), .Q(a_out[0]) );
  INVX3 U3 ( .A(rst), .Y(n1) );
endmodule


module top_DW01_inc_2 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
endmodule


module top_DW01_inc_3 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module top_DW01_inc_4 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module top_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [8:0] carry;

  ADDFXL U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADDFXL U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFXL U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFXL U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  INVXL U1 ( .A(B[0]), .Y(n8) );
  XNOR2XL U2 ( .A(A[5]), .B(carry[5]), .Y(DIFF[5]) );
  XNOR2XL U3 ( .A(A[6]), .B(carry[6]), .Y(DIFF[6]) );
  INVX1 U4 ( .A(B[2]), .Y(n6) );
  OR2X1 U5 ( .A(A[5]), .B(carry[5]), .Y(carry[6]) );
  CLKINVX1 U6 ( .A(B[4]), .Y(n4) );
  XNOR2X1 U7 ( .A(A[7]), .B(carry[7]), .Y(DIFF[7]) );
  NAND2X1 U8 ( .A(n2), .B(n3), .Y(carry[7]) );
  CLKINVX1 U9 ( .A(A[6]), .Y(n2) );
  CLKINVX1 U10 ( .A(carry[6]), .Y(n3) );
  CLKINVX1 U11 ( .A(B[3]), .Y(n5) );
  NAND2X1 U12 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U13 ( .A(B[1]), .Y(n7) );
  CLKINVX1 U14 ( .A(A[0]), .Y(n1) );
  XNOR2X1 U15 ( .A(n8), .B(A[0]), .Y(DIFF[0]) );
endmodule


module top ( clk, rst, start, m, n, k, done );
  input [3:0] m;
  input [3:0] n;
  input [3:0] k;
  input clk, rst, start;
  output done;
  wire   wr_en_out, load_en, \matrix_b[0][31] , \matrix_b[0][30] ,
         \matrix_b[0][29] , \matrix_b[0][28] , \matrix_b[0][27] ,
         \matrix_b[0][26] , \matrix_b[0][25] , \matrix_b[0][24] ,
         \matrix_b[0][23] , \matrix_b[0][22] , \matrix_b[0][21] ,
         \matrix_b[0][20] , \matrix_b[0][19] , \matrix_b[0][18] ,
         \matrix_b[0][17] , \matrix_b[0][16] , \matrix_b[0][15] ,
         \matrix_b[0][14] , \matrix_b[0][13] , \matrix_b[0][12] ,
         \matrix_b[0][11] , \matrix_b[0][10] , \matrix_b[0][9] ,
         \matrix_b[0][8] , \matrix_b[0][7] , \matrix_b[0][6] ,
         \matrix_b[0][5] , \matrix_b[0][4] , \matrix_b[0][3] ,
         \matrix_b[0][2] , \matrix_b[0][1] , \matrix_b[0][0] ,
         \matrix_b[1][15] , \matrix_b[1][14] , \matrix_b[1][13] ,
         \matrix_b[1][12] , \matrix_b[1][11] , \matrix_b[1][10] ,
         \matrix_b[1][9] , \matrix_b[1][8] , \matrix_b[1][7] ,
         \matrix_b[1][6] , \matrix_b[1][5] , \matrix_b[1][4] ,
         \matrix_b[1][3] , \matrix_b[1][2] , \matrix_b[1][1] ,
         \matrix_b[1][0] , \matrix_b[2][23] , \matrix_b[2][22] ,
         \matrix_b[2][21] , \matrix_b[2][20] , \matrix_b[2][19] ,
         \matrix_b[2][18] , \matrix_b[2][17] , \matrix_b[2][16] ,
         \matrix_b[2][15] , \matrix_b[2][14] , \matrix_b[2][13] ,
         \matrix_b[2][12] , \matrix_b[2][11] , \matrix_b[2][10] ,
         \matrix_b[2][9] , \matrix_b[2][8] , \matrix_b[3][31] ,
         \matrix_b[3][30] , \matrix_b[3][29] , \matrix_b[3][28] ,
         \matrix_b[3][27] , \matrix_b[3][26] , \matrix_b[3][25] ,
         \matrix_b[3][24] , \matrix_b[3][23] , \matrix_b[3][22] ,
         \matrix_b[3][21] , \matrix_b[3][20] , \matrix_b[3][19] ,
         \matrix_b[3][18] , \matrix_b[3][17] , \matrix_b[3][16] ,
         \matrix_b[4][31] , \matrix_b[4][30] , \matrix_b[4][29] ,
         \matrix_b[4][28] , \matrix_b[4][27] , \matrix_b[4][26] ,
         \matrix_b[4][25] , \matrix_b[4][24] , \matrix_b[4][7] ,
         \matrix_b[4][6] , \matrix_b[4][5] , \matrix_b[4][4] ,
         \matrix_b[4][3] , \matrix_b[4][2] , \matrix_b[4][1] ,
         \matrix_b[4][0] , \matrix_b[5][31] , \matrix_b[5][30] ,
         \matrix_b[5][29] , \matrix_b[5][28] , \matrix_b[5][27] ,
         \matrix_b[5][26] , \matrix_b[5][25] , \matrix_b[5][24] ,
         \matrix_b[5][15] , \matrix_b[5][14] , \matrix_b[5][13] ,
         \matrix_b[5][12] , \matrix_b[5][11] , \matrix_b[5][10] ,
         \matrix_b[5][9] , \matrix_b[5][8] , \matrix_b[5][7] ,
         \matrix_b[5][6] , \matrix_b[5][5] , \matrix_b[5][4] ,
         \matrix_b[5][3] , \matrix_b[5][2] , \matrix_b[5][1] ,
         \matrix_b[5][0] , \matrix_b[6][31] , \matrix_b[6][30] ,
         \matrix_b[6][29] , \matrix_b[6][28] , \matrix_b[6][27] ,
         \matrix_b[6][26] , \matrix_b[6][25] , \matrix_b[6][24] ,
         \matrix_b[6][23] , \matrix_b[6][22] , \matrix_b[6][21] ,
         \matrix_b[6][20] , \matrix_b[6][19] , \matrix_b[6][18] ,
         \matrix_b[6][17] , \matrix_b[6][16] , \matrix_b[6][15] ,
         \matrix_b[6][14] , \matrix_b[6][13] , \matrix_b[6][12] ,
         \matrix_b[6][11] , \matrix_b[6][10] , \matrix_b[6][9] ,
         \matrix_b[6][8] , \matrix_b[7][31] , \matrix_b[7][30] ,
         \matrix_b[7][29] , \matrix_b[7][28] , \matrix_b[7][27] ,
         \matrix_b[7][26] , \matrix_b[7][25] , \matrix_b[7][24] ,
         \matrix_b[7][23] , \matrix_b[7][22] , \matrix_b[7][21] ,
         \matrix_b[7][20] , \matrix_b[7][19] , \matrix_b[7][18] ,
         \matrix_b[7][17] , \matrix_b[7][16] , \matrix_b[8][31] ,
         \matrix_b[8][30] , \matrix_b[8][29] , \matrix_b[8][28] ,
         \matrix_b[8][27] , \matrix_b[8][26] , \matrix_b[8][25] ,
         \matrix_b[8][24] , \matrix_b[8][23] , \matrix_b[8][22] ,
         \matrix_b[8][21] , \matrix_b[8][20] , \matrix_b[8][19] ,
         \matrix_b[8][18] , \matrix_b[8][17] , \matrix_b[8][16] ,
         \matrix_b[8][15] , \matrix_b[8][14] , \matrix_b[8][13] ,
         \matrix_b[8][12] , \matrix_b[8][11] , \matrix_b[8][10] ,
         \matrix_b[8][9] , \matrix_b[8][8] , \matrix_b[8][7] ,
         \matrix_b[8][6] , \matrix_b[8][5] , \matrix_b[8][4] ,
         \matrix_b[8][3] , \matrix_b[8][2] , \matrix_b[8][1] ,
         \matrix_b[8][0] , N241, N243, N244, N247, N252, N253, N254, N257,
         N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268,
         N269, N270, N271, N272, N630, N631, N632, N633, N634, N635, N636,
         N637, N638, N639, N640, N712, N713, N714, N715, N719, N720, N721,
         N722, N726, N727, N731, N732, N733, N780, N781, N782, N783, N784,
         N785, N786, N787, N788, N789, N791, N793, N802, N803, N804, N805,
         N806, N807, N808, N809, N892, N894, N896, N898, N912, n163, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n629,
         n630, n631, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n779, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n822, n823, n825, n827, n828, n829, n831, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1146,
         n1151, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1272, n1274, n1275, n1276, n1277, n1278,
         n1279, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, N798,
         N797, N796, N795, N794, \add_357/carry[3] , \add_357/carry[2] ,
         \add_332_3/carry[2] , \add_332/carry[3] , \add_332/carry[2] ,
         \add_331/carry[3] , \add_331/carry[2] , \sub_142/carry[4] ,
         \add_357_2/carry[4] , \add_357_2/carry[3] ,
         \add_1_root_sub_0_root_sub_359_2/carry[3] ,
         \add_1_root_sub_0_root_sub_359_2/carry[2] , n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912;
  wire   [7:0] index_a;
  wire   [31:0] data_in_a;
  wire   [31:0] data_out_a;
  wire   [7:0] index_b;
  wire   [31:0] data_in_b;
  wire   [31:0] data_out_b;
  wire   [7:0] index_out;
  wire   [31:0] data_in_o;
  wire   [1:0] cur_state;
  wire   [1:0] next_state;
  wire   [5:0] l;
  wire   [10:0] counter;
  wire   [7:0] a11;
  wire   [7:0] a12;
  wire   [7:0] a13;
  wire   [7:0] a14;
  wire   [7:0] b11;
  wire   [7:0] b12;
  wire   [7:0] b21;
  wire   [7:0] b13;
  wire   [7:0] b22;
  wire   [7:0] b31;
  wire   [7:0] b14;
  wire   [7:0] b23;
  wire   [7:0] b32;
  wire   [7:0] b41;
  wire   [7:0] b24;
  wire   [7:0] b33;
  wire   [7:0] b42;
  wire   [7:0] b34;
  wire   [7:0] b43;
  wire   [7:0] b44;
  wire   [7:0] w11;
  wire   [7:0] w21;
  wire   [7:0] w31;
  wire   [7:0] w41;
  wire   [7:0] w12;
  wire   [7:0] w22;
  wire   [7:0] w32;
  wire   [7:0] w42;
  wire   [7:0] w13;
  wire   [7:0] w23;
  wire   [7:0] w33;
  wire   [7:0] w43;
  wire   [7:0] w14;
  wire   [7:0] w24;
  wire   [7:0] w34;
  wire   [7:0] w44;
  wire   [23:0] temp1;
  wire   [7:0] psum1;
  wire   [7:0] psum2;
  wire   [7:0] psum3;
  wire   [7:0] psum4;
  wire   [7:0] a21;
  wire   [7:0] a22;
  wire   [7:0] a23;
  wire   [7:0] a24;
  wire   [7:0] a31;
  wire   [7:0] a32;
  wire   [7:0] a33;
  wire   [7:0] a34;
  wire   [7:0] a41;
  wire   [7:0] a42;
  wire   [7:0] a43;
  wire   [7:0] a44;
  assign done = 1'b1;
  assign N241 = k[1];
  assign N247 = k[2];
  assign N785 = k[0];

  global_buffer_0 GBUFF_A ( .clk(clk), .rst(n1521), .wr_en(1'b0), .index({
        index_a[7:5], n1695, n1694, index_a[2], n1691, n1689}), .data_in({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_out(data_out_a) );
  global_buffer_2 GBUFF_B ( .clk(clk), .rst(n1521), .wr_en(1'b0), .index({
        index_b[7:5], n1688, n1687, n1685, n1683, n1681}), .data_in({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_out(data_out_b) );
  global_buffer_1 GBUFF_OUT ( .clk(clk), .rst(n1521), .wr_en(wr_en_out), 
        .index(index_out), .data_in(data_in_o) );
  pe_0 pe_w11 ( .clk(clk), .rst(n1521), .a(a11), .b(b11), .psum(psum1), 
        .a_out(a21), .out(w11) );
  pe_15 pe_w12 ( .clk(clk), .rst(n1521), .a(a12), .b(b12), .psum(w11), .a_out(
        a22), .out(w12) );
  pe_14 pe_w13 ( .clk(clk), .rst(n1521), .a(a13), .b(b13), .psum(w12), .a_out(
        a23), .out(w13) );
  pe_13 pe_w14 ( .clk(clk), .rst(n1521), .a(a14), .b(b14), .psum(w13), .a_out(
        a24), .out(w14) );
  pe_12 pe_w21 ( .clk(clk), .rst(n1521), .a(a21), .b(b21), .psum(psum2), 
        .a_out(a31), .out(w21) );
  pe_11 pe_w22 ( .clk(clk), .rst(n1521), .a(a22), .b(b22), .psum(w21), .a_out(
        a32), .out(w22) );
  pe_10 pe_w23 ( .clk(clk), .rst(n1521), .a(a23), .b(b23), .psum(w22), .a_out(
        a33), .out(w23) );
  pe_9 pe_w24 ( .clk(clk), .rst(n1521), .a(a24), .b(b24), .psum(w23), .a_out(
        a34), .out(w24) );
  pe_8 pe_w31 ( .clk(clk), .rst(n1521), .a(a31), .b(b31), .psum(psum3), 
        .a_out(a41), .out(w31) );
  pe_7 pe_w32 ( .clk(clk), .rst(n1521), .a(a32), .b(b32), .psum(w31), .a_out(
        a42), .out(w32) );
  pe_6 pe_w33 ( .clk(clk), .rst(n1521), .a(a33), .b(b33), .psum(w32), .a_out(
        a43), .out(w33) );
  pe_5 pe_w34 ( .clk(clk), .rst(n1521), .a(a34), .b(b34), .psum(w33), .a_out(
        a44), .out(w34) );
  pe_4 pe_w41 ( .clk(clk), .rst(n1521), .a(a41), .b(b41), .psum(psum4), .out(
        w41) );
  pe_3 pe_w42 ( .clk(clk), .rst(n1521), .a(a42), .b(b42), .psum(w41), .out(w42) );
  pe_2 pe_w43 ( .clk(clk), .rst(n1521), .a(a43), .b(b43), .psum(w42), .out(w43) );
  pe_1 pe_w44 ( .clk(clk), .rst(n1521), .a(a44), .b(b44), .psum(w43), .out(w44) );
  top_DW01_inc_2 add_289 ( .A({n1621, n1622, n1623, n1624, n1625, n1626, n1627, 
        n1628, n1629, n1630, n1631}), .SUM({N640, N639, N638, N637, N636, N635, 
        N634, N633, N632, N631, N630}) );
  top_DW01_inc_3 add_151 ( .A({index_b[7:5], n1688, n1687, n1685, n1683, n1681}), .SUM({N272, N271, N270, N269, N268, N267, N266, N265}) );
  top_DW01_inc_4 add_150 ( .A({index_a[7:5], n1695, n1694, index_a[2], n1691, 
        n1689}), .SUM({N264, N263, N262, N261, N260, N259, N258, N257}) );
  top_DW01_sub_2 sub_0_root_sub_0_root_sub_359_2 ( .A({n1624, n1625, n1626, 
        n1627, n1628, n1629, n1630, n1631}), .B({1'b0, 1'b0, 1'b0, N798, N797, 
        N796, N795, N794}), .CI(1'b0), .DIFF({N809, N808, N807, N806, N805, 
        N804, N803, N802}) );
  EDFFX1 \matrix_b_reg[6][7]  ( .D(data_out_b[7]), .E(n1556), .CK(clk), .QN(
        n586) );
  EDFFX1 \matrix_b_reg[6][6]  ( .D(data_out_b[6]), .E(n1556), .CK(clk), .QN(
        n587) );
  EDFFX1 \matrix_b_reg[6][5]  ( .D(data_out_b[5]), .E(n1556), .CK(clk), .QN(
        n588) );
  EDFFX1 \matrix_b_reg[6][4]  ( .D(data_out_b[4]), .E(n1556), .CK(clk), .QN(
        n589) );
  EDFFX1 \matrix_b_reg[6][3]  ( .D(data_out_b[3]), .E(n1556), .CK(clk), .QN(
        n590) );
  EDFFX1 \matrix_b_reg[6][2]  ( .D(data_out_b[2]), .E(n1556), .CK(clk), .QN(
        n591) );
  EDFFX1 \matrix_b_reg[6][1]  ( .D(data_out_b[1]), .E(n1556), .CK(clk), .QN(
        n592) );
  EDFFX1 \matrix_b_reg[6][0]  ( .D(data_out_b[0]), .E(n1556), .CK(clk), .QN(
        n593) );
  EDFFX1 \temp3_reg[0]  ( .D(n954), .E(n1562), .CK(clk), .QN(n708) );
  EDFFX1 \temp3_reg[1]  ( .D(n938), .E(n1562), .CK(clk), .QN(n707) );
  EDFFX1 \temp3_reg[2]  ( .D(n935), .E(n1632), .CK(clk), .QN(n706) );
  EDFFX1 \temp3_reg[3]  ( .D(n932), .E(n1632), .CK(clk), .QN(n705) );
  EDFFX1 \temp3_reg[4]  ( .D(n929), .E(n1632), .CK(clk), .QN(n704) );
  EDFFX1 \temp3_reg[5]  ( .D(n926), .E(n1632), .CK(clk), .QN(n703) );
  EDFFX1 \temp3_reg[6]  ( .D(n923), .E(n1632), .CK(clk), .QN(n702) );
  EDFFX1 \temp3_reg[7]  ( .D(n920), .E(n1632), .CK(clk), .QN(n701) );
  EDFFX1 \temp2_reg[8]  ( .D(n900), .E(n1562), .CK(clk), .QN(n732) );
  EDFFX1 \temp2_reg[9]  ( .D(n897), .E(n1562), .CK(clk), .QN(n731) );
  EDFFX1 \temp2_reg[10]  ( .D(n894), .E(n1632), .CK(clk), .QN(n730) );
  EDFFX1 \temp2_reg[11]  ( .D(n891), .E(n1632), .CK(clk), .QN(n729) );
  EDFFX1 \temp2_reg[12]  ( .D(n888), .E(n1632), .CK(clk), .QN(n728) );
  EDFFX1 \temp2_reg[13]  ( .D(n885), .E(n1632), .CK(clk), .QN(n727) );
  EDFFX1 \temp2_reg[14]  ( .D(n882), .E(n1632), .CK(clk), .QN(n726) );
  EDFFX1 \temp2_reg[15]  ( .D(n879), .E(n1632), .CK(clk), .QN(n725) );
  EDFFTRX1 work_fin_reg ( .RN(n1906), .D(1'b1), .E(n1555), .CK(clk), .QN(n741)
         );
  EDFFX1 \temp1_reg[16]  ( .D(n823), .E(n1632), .CK(clk), .Q(temp1[16]) );
  EDFFX1 \temp1_reg[17]  ( .D(n825), .E(n1632), .CK(clk), .Q(temp1[17]) );
  EDFFX1 \temp1_reg[18]  ( .D(n827), .E(n1632), .CK(clk), .Q(temp1[18]) );
  EDFFX1 \temp1_reg[19]  ( .D(n829), .E(n1632), .CK(clk), .Q(temp1[19]) );
  EDFFX1 \temp1_reg[20]  ( .D(n831), .E(n1632), .CK(clk), .Q(temp1[20]) );
  EDFFX1 \temp1_reg[21]  ( .D(n833), .E(n1632), .CK(clk), .Q(temp1[21]) );
  EDFFX1 \temp1_reg[22]  ( .D(n835), .E(n1632), .CK(clk), .Q(temp1[22]) );
  EDFFX1 \temp1_reg[23]  ( .D(n837), .E(n1632), .CK(clk), .Q(temp1[23]) );
  EDFFX1 \matrix_b_reg[6][15]  ( .D(data_out_b[15]), .E(n1633), .CK(clk), .Q(
        \matrix_b[6][15] ) );
  EDFFX1 \matrix_b_reg[6][14]  ( .D(data_out_b[14]), .E(n1633), .CK(clk), .Q(
        \matrix_b[6][14] ) );
  EDFFX1 \matrix_b_reg[6][13]  ( .D(data_out_b[13]), .E(n1633), .CK(clk), .Q(
        \matrix_b[6][13] ) );
  EDFFX1 \matrix_b_reg[6][12]  ( .D(data_out_b[12]), .E(n1633), .CK(clk), .Q(
        \matrix_b[6][12] ) );
  EDFFX1 \matrix_b_reg[6][11]  ( .D(data_out_b[11]), .E(n1633), .CK(clk), .Q(
        \matrix_b[6][11] ) );
  EDFFX1 \matrix_b_reg[6][10]  ( .D(data_out_b[10]), .E(n1633), .CK(clk), .Q(
        \matrix_b[6][10] ) );
  EDFFX1 \matrix_b_reg[6][9]  ( .D(data_out_b[9]), .E(n1633), .CK(clk), .Q(
        \matrix_b[6][9] ) );
  EDFFX1 \matrix_b_reg[6][8]  ( .D(data_out_b[8]), .E(n1633), .CK(clk), .Q(
        \matrix_b[6][8] ) );
  EDFFX1 \matrix_a_reg[1][23]  ( .D(n1593), .E(n1568), .CK(clk), .QN(n266) );
  EDFFX1 \matrix_a_reg[1][22]  ( .D(n1592), .E(n1568), .CK(clk), .QN(n267) );
  EDFFX1 \matrix_a_reg[1][21]  ( .D(n1591), .E(n1568), .CK(clk), .QN(n268) );
  EDFFX1 \matrix_a_reg[1][20]  ( .D(n1590), .E(n1636), .CK(clk), .QN(n269) );
  EDFFX1 \matrix_a_reg[1][19]  ( .D(n1589), .E(n1636), .CK(clk), .QN(n270) );
  EDFFX1 \matrix_a_reg[1][18]  ( .D(n1588), .E(n1636), .CK(clk), .QN(n271) );
  EDFFX1 \matrix_a_reg[1][17]  ( .D(n1587), .E(n1636), .CK(clk), .QN(n272) );
  EDFFX1 \matrix_a_reg[1][16]  ( .D(n1586), .E(n1636), .CK(clk), .QN(n273) );
  EDFFX1 \matrix_a_reg[6][23]  ( .D(n1593), .E(n1557), .CK(clk), .QN(n426) );
  EDFFX1 \matrix_a_reg[6][22]  ( .D(n1592), .E(n1557), .CK(clk), .QN(n427) );
  EDFFX1 \matrix_a_reg[6][21]  ( .D(n1591), .E(n1557), .CK(clk), .QN(n428) );
  EDFFX1 \matrix_a_reg[6][20]  ( .D(n1590), .E(n1557), .CK(clk), .QN(n429) );
  EDFFX1 \matrix_a_reg[6][19]  ( .D(n1589), .E(n1557), .CK(clk), .QN(n430) );
  EDFFX1 \matrix_a_reg[6][18]  ( .D(n1588), .E(n1557), .CK(clk), .QN(n431) );
  EDFFX1 \matrix_a_reg[6][17]  ( .D(n1587), .E(n1557), .CK(clk), .QN(n432) );
  EDFFX1 \matrix_a_reg[6][16]  ( .D(n1586), .E(n1557), .CK(clk), .QN(n433) );
  EDFFX1 \matrix_a_reg[6][7]  ( .D(data_out_a[7]), .E(n1635), .CK(clk), .QN(
        n442) );
  EDFFX1 \matrix_a_reg[6][6]  ( .D(data_out_a[6]), .E(n1635), .CK(clk), .QN(
        n443) );
  EDFFX1 \matrix_a_reg[6][5]  ( .D(data_out_a[5]), .E(n1635), .CK(clk), .QN(
        n444) );
  EDFFX1 \matrix_a_reg[6][4]  ( .D(data_out_a[4]), .E(n1635), .CK(clk), .QN(
        n445) );
  EDFFX1 \matrix_a_reg[6][3]  ( .D(data_out_a[3]), .E(n1635), .CK(clk), .QN(
        n446) );
  EDFFX1 \matrix_a_reg[6][2]  ( .D(data_out_a[2]), .E(n1635), .CK(clk), .QN(
        n447) );
  EDFFX1 \matrix_a_reg[6][1]  ( .D(data_out_a[1]), .E(n1635), .CK(clk), .QN(
        n448) );
  EDFFX1 \matrix_a_reg[6][0]  ( .D(data_out_a[0]), .E(n1635), .CK(clk), .QN(
        n449) );
  DFFX1 \matrix_b_reg[3][15]  ( .D(n1467), .CK(clk), .QN(n546) );
  DFFX1 \matrix_b_reg[3][14]  ( .D(n1468), .CK(clk), .QN(n547) );
  DFFX1 \matrix_b_reg[3][13]  ( .D(n1469), .CK(clk), .QN(n548) );
  DFFX1 \matrix_b_reg[3][12]  ( .D(n1470), .CK(clk), .QN(n549) );
  DFFX1 \matrix_b_reg[3][11]  ( .D(n1471), .CK(clk), .QN(n550) );
  DFFX1 \matrix_b_reg[3][10]  ( .D(n1472), .CK(clk), .QN(n551) );
  DFFX1 \matrix_b_reg[3][9]  ( .D(n1473), .CK(clk), .QN(n552) );
  DFFX1 \matrix_b_reg[3][8]  ( .D(n1474), .CK(clk), .QN(n553) );
  DFFX1 \matrix_b_reg[3][7]  ( .D(n1483), .CK(clk), .QN(n554) );
  DFFX1 \matrix_b_reg[3][6]  ( .D(n1484), .CK(clk), .QN(n555) );
  DFFX1 \matrix_b_reg[3][5]  ( .D(n1485), .CK(clk), .QN(n556) );
  DFFX1 \matrix_b_reg[3][4]  ( .D(n1486), .CK(clk), .QN(n557) );
  DFFX1 \matrix_b_reg[3][3]  ( .D(n1487), .CK(clk), .QN(n558) );
  DFFX1 \matrix_b_reg[3][2]  ( .D(n1488), .CK(clk), .QN(n559) );
  DFFX1 \matrix_b_reg[3][1]  ( .D(n1489), .CK(clk), .QN(n560) );
  DFFX1 \matrix_b_reg[3][0]  ( .D(n1490), .CK(clk), .QN(n561) );
  DFFQX1 load_en_reg ( .D(n1507), .CK(clk), .Q(load_en) );
  EDFFX1 \matrix_a_reg[6][31]  ( .D(data_out_a[31]), .E(n1635), .CK(clk), .QN(
        n418) );
  EDFFX1 \matrix_a_reg[6][30]  ( .D(data_out_a[30]), .E(n1635), .CK(clk), .QN(
        n419) );
  EDFFX1 \matrix_a_reg[6][29]  ( .D(data_out_a[29]), .E(n1635), .CK(clk), .QN(
        n420) );
  EDFFX1 \matrix_a_reg[6][28]  ( .D(data_out_a[28]), .E(n1635), .CK(clk), .QN(
        n421) );
  EDFFX1 \matrix_a_reg[6][27]  ( .D(data_out_a[27]), .E(n1635), .CK(clk), .QN(
        n422) );
  EDFFX1 \matrix_a_reg[6][26]  ( .D(data_out_a[26]), .E(n1635), .CK(clk), .QN(
        n423) );
  EDFFX1 \matrix_a_reg[6][25]  ( .D(data_out_a[25]), .E(n1557), .CK(clk), .QN(
        n424) );
  EDFFX1 \matrix_a_reg[6][24]  ( .D(data_out_a[24]), .E(n1557), .CK(clk), .QN(
        n425) );
  EDFFX1 \matrix_a_reg[6][15]  ( .D(n1585), .E(n1557), .CK(clk), .QN(n434) );
  EDFFX1 \matrix_a_reg[6][14]  ( .D(n1584), .E(n1557), .CK(clk), .QN(n435) );
  EDFFX1 \matrix_a_reg[6][13]  ( .D(n1583), .E(n1635), .CK(clk), .QN(n436) );
  EDFFX1 \matrix_a_reg[6][12]  ( .D(n1582), .E(n1635), .CK(clk), .QN(n437) );
  EDFFX1 \matrix_a_reg[6][11]  ( .D(n1581), .E(n1635), .CK(clk), .QN(n438) );
  EDFFX1 \matrix_a_reg[6][10]  ( .D(n1580), .E(n1635), .CK(clk), .QN(n439) );
  EDFFX1 \matrix_a_reg[6][9]  ( .D(n1579), .E(n1635), .CK(clk), .QN(n440) );
  EDFFX1 \matrix_a_reg[6][8]  ( .D(n1578), .E(n1635), .CK(clk), .QN(n441) );
  EDFFX1 \matrix_a_reg[1][15]  ( .D(n1585), .E(n1636), .CK(clk), .QN(n274) );
  EDFFX1 \matrix_a_reg[1][14]  ( .D(n1584), .E(n1636), .CK(clk), .QN(n275) );
  EDFFX1 \matrix_a_reg[1][13]  ( .D(n1583), .E(n1636), .CK(clk), .QN(n276) );
  EDFFX1 \matrix_a_reg[1][12]  ( .D(n1582), .E(n1636), .CK(clk), .QN(n277) );
  EDFFX1 \matrix_a_reg[1][11]  ( .D(n1581), .E(n1636), .CK(clk), .QN(n278) );
  EDFFX1 \matrix_a_reg[1][10]  ( .D(n1580), .E(n1636), .CK(clk), .QN(n279) );
  EDFFX1 \matrix_a_reg[1][9]  ( .D(n1579), .E(n1636), .CK(clk), .QN(n280) );
  EDFFX1 \matrix_a_reg[1][8]  ( .D(n1578), .E(n1636), .CK(clk), .QN(n281) );
  EDFFX1 \index_out_reg[4]  ( .D(N806), .E(n1680), .CK(clk), .Q(index_out[4])
         );
  EDFFX1 \index_out_reg[2]  ( .D(N804), .E(n1680), .CK(clk), .Q(index_out[2])
         );
  DFFX1 \matrix_a_reg[3][23]  ( .D(n1371), .CK(clk), .QN(n330) );
  DFFX1 \matrix_a_reg[3][22]  ( .D(n1372), .CK(clk), .QN(n331) );
  DFFX1 \matrix_a_reg[3][21]  ( .D(n1373), .CK(clk), .QN(n332) );
  DFFX1 \matrix_a_reg[3][20]  ( .D(n1374), .CK(clk), .QN(n333) );
  DFFX1 \matrix_a_reg[3][19]  ( .D(n1375), .CK(clk), .QN(n334) );
  DFFX1 \matrix_a_reg[3][18]  ( .D(n1376), .CK(clk), .QN(n335) );
  DFFX1 \matrix_a_reg[3][17]  ( .D(n1377), .CK(clk), .QN(n336) );
  DFFX1 \matrix_a_reg[3][16]  ( .D(n1378), .CK(clk), .QN(n337) );
  DFFX1 \matrix_a_reg[3][7]  ( .D(n1387), .CK(clk), .QN(n346) );
  DFFX1 \matrix_a_reg[3][6]  ( .D(n1388), .CK(clk), .QN(n347) );
  DFFX1 \matrix_a_reg[3][5]  ( .D(n1389), .CK(clk), .QN(n348) );
  DFFX1 \matrix_a_reg[3][4]  ( .D(n1390), .CK(clk), .QN(n349) );
  DFFX1 \matrix_a_reg[3][3]  ( .D(n1391), .CK(clk), .QN(n350) );
  DFFX1 \matrix_a_reg[3][2]  ( .D(n1392), .CK(clk), .QN(n351) );
  DFFX1 \matrix_a_reg[3][1]  ( .D(n1393), .CK(clk), .QN(n352) );
  DFFX1 \matrix_a_reg[3][0]  ( .D(n1394), .CK(clk), .QN(n353) );
  DFFX1 \matrix_a_reg[3][31]  ( .D(n1363), .CK(clk), .QN(n322) );
  DFFX1 \matrix_a_reg[3][30]  ( .D(n1364), .CK(clk), .QN(n323) );
  DFFX1 \matrix_a_reg[3][29]  ( .D(n1365), .CK(clk), .QN(n324) );
  DFFX1 \matrix_a_reg[3][28]  ( .D(n1366), .CK(clk), .QN(n325) );
  DFFX1 \matrix_a_reg[3][27]  ( .D(n1367), .CK(clk), .QN(n326) );
  DFFX1 \matrix_a_reg[3][26]  ( .D(n1368), .CK(clk), .QN(n327) );
  DFFX1 \matrix_a_reg[3][25]  ( .D(n1369), .CK(clk), .QN(n328) );
  DFFX1 \matrix_a_reg[3][24]  ( .D(n1370), .CK(clk), .QN(n329) );
  DFFX1 \matrix_a_reg[3][15]  ( .D(n1379), .CK(clk), .QN(n338) );
  DFFX1 \matrix_a_reg[3][14]  ( .D(n1380), .CK(clk), .QN(n339) );
  DFFX1 \matrix_a_reg[3][13]  ( .D(n1381), .CK(clk), .QN(n340) );
  DFFX1 \matrix_a_reg[3][12]  ( .D(n1382), .CK(clk), .QN(n341) );
  DFFX1 \matrix_a_reg[3][11]  ( .D(n1383), .CK(clk), .QN(n342) );
  DFFX1 \matrix_a_reg[3][10]  ( .D(n1384), .CK(clk), .QN(n343) );
  DFFX1 \matrix_a_reg[3][9]  ( .D(n1385), .CK(clk), .QN(n344) );
  DFFX1 \matrix_a_reg[3][8]  ( .D(n1386), .CK(clk), .QN(n345) );
  DFFQX1 \index_a_reg[2]  ( .D(n1504), .CK(clk), .Q(index_a[2]) );
  DFFX1 \b43_reg[7]  ( .D(n1451), .CK(clk), .Q(b43[7]), .QN(n667) );
  DFFX1 \b44_reg[7]  ( .D(n1475), .CK(clk), .Q(b44[7]), .QN(n675) );
  DFFX1 \b12_reg[7]  ( .D(n1427), .CK(clk), .Q(b12[7]), .QN(n635) );
  DFFX1 \b13_reg[7]  ( .D(n1443), .CK(clk), .Q(b13[7]), .QN(n651) );
  DFFX1 \b22_reg[7]  ( .D(n1435), .CK(clk), .Q(b22[7]), .QN(n643) );
  DFFX1 \b34_reg[7]  ( .D(n1459), .CK(clk), .Q(b34[7]), .QN(n659) );
  EDFFX1 \index_out_reg[5]  ( .D(N807), .E(n1680), .CK(clk), .Q(index_out[5])
         );
  DFFQX1 \b41_reg[7]  ( .D(n1419), .CK(clk), .Q(b41[7]) );
  DFFQX1 \b11_reg[7]  ( .D(n1395), .CK(clk), .Q(b11[7]) );
  DFFQX1 \b21_reg[7]  ( .D(n1403), .CK(clk), .Q(b21[7]) );
  DFFQX1 \b31_reg[7]  ( .D(n1411), .CK(clk), .Q(b31[7]) );
  EDFFX1 \l_reg[4]  ( .D(N254), .E(n1907), .CK(clk), .Q(l[4]) );
  EDFFX1 \l_reg[3]  ( .D(N253), .E(n1907), .CK(clk), .Q(l[3]) );
  DFFQX1 \b42_reg[7]  ( .D(n1881), .CK(clk), .Q(b42[7]) );
  DFFQX1 \b14_reg[7]  ( .D(n1889), .CK(clk), .Q(b14[7]) );
  DFFQX1 \b23_reg[7]  ( .D(n1897), .CK(clk), .Q(b23[7]) );
  DFFQX1 \b24_reg[7]  ( .D(n1865), .CK(clk), .Q(b24[7]) );
  DFFQX1 \b32_reg[7]  ( .D(n1905), .CK(clk), .Q(b32[7]) );
  DFFQX1 \b33_reg[7]  ( .D(n1873), .CK(clk), .Q(b33[7]) );
  EDFFX1 \l_reg[5]  ( .D(N254), .E(n1907), .CK(clk), .Q(l[5]) );
  DFFQX1 \index_b_reg[3]  ( .D(n1494), .CK(clk), .Q(index_b[3]) );
  DFFQX1 \index_b_reg[4]  ( .D(n1493), .CK(clk), .Q(index_b[4]) );
  DFFQX1 \index_a_reg[3]  ( .D(n1503), .CK(clk), .Q(index_a[3]) );
  DFFQX1 \index_a_reg[4]  ( .D(n1502), .CK(clk), .Q(index_a[4]) );
  DFFQX1 \a14_reg[7]  ( .D(n1355), .CK(clk), .Q(a14[7]) );
  DFFQX1 \a11_reg[7]  ( .D(n1331), .CK(clk), .Q(a11[7]) );
  DFFQX1 \a12_reg[7]  ( .D(n1339), .CK(clk), .Q(a12[7]) );
  DFFQX1 \a13_reg[7]  ( .D(n1347), .CK(clk), .Q(a13[7]) );
  DFFRX1 \cur_state_reg[0]  ( .D(next_state[0]), .CK(clk), .RN(n1851), .Q(
        cur_state[0]), .QN(n225) );
  DFFQX1 \index_b_reg[0]  ( .D(n1497), .CK(clk), .Q(index_b[0]) );
  DFFQX1 \index_b_reg[1]  ( .D(n1496), .CK(clk), .Q(index_b[1]) );
  DFFQX1 \index_b_reg[2]  ( .D(n1495), .CK(clk), .Q(index_b[2]) );
  DFFQX1 \index_a_reg[0]  ( .D(n1506), .CK(clk), .Q(index_a[0]) );
  DFFQX1 \index_a_reg[1]  ( .D(n1505), .CK(clk), .Q(index_a[1]) );
  EDFFX1 \index_out_reg[3]  ( .D(N805), .E(n1680), .CK(clk), .Q(index_out[3])
         );
  EDFFX1 \index_out_reg[1]  ( .D(N803), .E(n1680), .CK(clk), .Q(index_out[1])
         );
  EDFFX1 \index_out_reg[0]  ( .D(N802), .E(n1680), .CK(clk), .Q(index_out[0])
         );
  DFFQX1 \index_a_reg[7]  ( .D(n1508), .CK(clk), .Q(index_a[7]) );
  DFFQX1 \index_b_reg[7]  ( .D(n1498), .CK(clk), .Q(index_b[7]) );
  DFFRX1 \cur_state_reg[1]  ( .D(next_state[1]), .CK(clk), .RN(n1851), .Q(
        cur_state[1]), .QN(n163) );
  DFFX1 \b43_reg[6]  ( .D(n1452), .CK(clk), .Q(b43[6]), .QN(n668) );
  DFFX1 \b44_reg[6]  ( .D(n1476), .CK(clk), .Q(b44[6]), .QN(n676) );
  DFFX1 \b12_reg[6]  ( .D(n1428), .CK(clk), .Q(b12[6]), .QN(n636) );
  DFFX1 \b13_reg[6]  ( .D(n1444), .CK(clk), .Q(b13[6]), .QN(n652) );
  DFFX1 \b22_reg[6]  ( .D(n1436), .CK(clk), .Q(b22[6]), .QN(n644) );
  DFFX1 \b34_reg[6]  ( .D(n1460), .CK(clk), .Q(b34[6]), .QN(n660) );
  DFFX1 \b43_reg[5]  ( .D(n1453), .CK(clk), .Q(b43[5]), .QN(n669) );
  DFFX1 \b43_reg[4]  ( .D(n1454), .CK(clk), .Q(b43[4]), .QN(n670) );
  DFFX1 \b44_reg[5]  ( .D(n1477), .CK(clk), .Q(b44[5]), .QN(n677) );
  DFFX1 \b44_reg[4]  ( .D(n1478), .CK(clk), .Q(b44[4]), .QN(n678) );
  DFFX1 \b12_reg[5]  ( .D(n1429), .CK(clk), .Q(b12[5]), .QN(n637) );
  DFFX1 \b12_reg[4]  ( .D(n1430), .CK(clk), .Q(b12[4]), .QN(n638) );
  DFFX1 \b13_reg[5]  ( .D(n1445), .CK(clk), .Q(b13[5]), .QN(n653) );
  DFFX1 \b13_reg[4]  ( .D(n1446), .CK(clk), .Q(b13[4]), .QN(n654) );
  DFFX1 \b22_reg[5]  ( .D(n1437), .CK(clk), .Q(b22[5]), .QN(n645) );
  DFFX1 \b22_reg[4]  ( .D(n1438), .CK(clk), .Q(b22[4]), .QN(n646) );
  DFFX1 \b34_reg[5]  ( .D(n1461), .CK(clk), .Q(b34[5]), .QN(n661) );
  DFFX1 \b34_reg[4]  ( .D(n1462), .CK(clk), .Q(b34[4]), .QN(n662) );
  DFFQX1 \b41_reg[6]  ( .D(n1420), .CK(clk), .Q(b41[6]) );
  DFFQX1 \b11_reg[6]  ( .D(n1396), .CK(clk), .Q(b11[6]) );
  DFFQX1 \b21_reg[6]  ( .D(n1404), .CK(clk), .Q(b21[6]) );
  DFFQX1 \b31_reg[6]  ( .D(n1412), .CK(clk), .Q(b31[6]) );
  DFFQX1 \b42_reg[6]  ( .D(n1880), .CK(clk), .Q(b42[6]) );
  DFFQX1 \b14_reg[6]  ( .D(n1888), .CK(clk), .Q(b14[6]) );
  DFFQX1 \b23_reg[6]  ( .D(n1896), .CK(clk), .Q(b23[6]) );
  DFFQX1 \b24_reg[6]  ( .D(n1864), .CK(clk), .Q(b24[6]) );
  DFFQX1 \b32_reg[6]  ( .D(n1904), .CK(clk), .Q(b32[6]) );
  DFFQX1 \b33_reg[6]  ( .D(n1872), .CK(clk), .Q(b33[6]) );
  DFFQX1 \b41_reg[5]  ( .D(n1421), .CK(clk), .Q(b41[5]) );
  DFFQX1 \b41_reg[4]  ( .D(n1422), .CK(clk), .Q(b41[4]) );
  DFFQX1 \b11_reg[5]  ( .D(n1397), .CK(clk), .Q(b11[5]) );
  DFFQX1 \b11_reg[4]  ( .D(n1398), .CK(clk), .Q(b11[4]) );
  DFFQX1 \b21_reg[5]  ( .D(n1405), .CK(clk), .Q(b21[5]) );
  DFFQX1 \b21_reg[4]  ( .D(n1406), .CK(clk), .Q(b21[4]) );
  DFFQX1 \b31_reg[5]  ( .D(n1413), .CK(clk), .Q(b31[5]) );
  DFFQX1 \b31_reg[4]  ( .D(n1414), .CK(clk), .Q(b31[4]) );
  DFFQX1 \b42_reg[5]  ( .D(n1879), .CK(clk), .Q(b42[5]) );
  DFFQX1 \b42_reg[4]  ( .D(n1878), .CK(clk), .Q(b42[4]) );
  DFFQX1 \b14_reg[5]  ( .D(n1887), .CK(clk), .Q(b14[5]) );
  DFFQX1 \b14_reg[4]  ( .D(n1886), .CK(clk), .Q(b14[4]) );
  DFFQX1 \b23_reg[5]  ( .D(n1895), .CK(clk), .Q(b23[5]) );
  DFFQX1 \b23_reg[4]  ( .D(n1894), .CK(clk), .Q(b23[4]) );
  DFFQX1 \b24_reg[5]  ( .D(n1863), .CK(clk), .Q(b24[5]) );
  DFFQX1 \b24_reg[4]  ( .D(n1862), .CK(clk), .Q(b24[4]) );
  DFFQX1 \b32_reg[5]  ( .D(n1903), .CK(clk), .Q(b32[5]) );
  DFFQX1 \b32_reg[4]  ( .D(n1902), .CK(clk), .Q(b32[4]) );
  DFFQX1 \b33_reg[5]  ( .D(n1871), .CK(clk), .Q(b33[5]) );
  DFFQX1 \b33_reg[4]  ( .D(n1870), .CK(clk), .Q(b33[4]) );
  DFFQX1 \a14_reg[6]  ( .D(n1356), .CK(clk), .Q(a14[6]) );
  DFFQX1 \a11_reg[6]  ( .D(n1332), .CK(clk), .Q(a11[6]) );
  DFFQX1 \a12_reg[6]  ( .D(n1340), .CK(clk), .Q(a12[6]) );
  DFFQX1 \a13_reg[6]  ( .D(n1348), .CK(clk), .Q(a13[6]) );
  DFFQX1 \a14_reg[5]  ( .D(n1357), .CK(clk), .Q(a14[5]) );
  DFFQX1 \a14_reg[4]  ( .D(n1358), .CK(clk), .Q(a14[4]) );
  DFFQX1 \a11_reg[5]  ( .D(n1333), .CK(clk), .Q(a11[5]) );
  DFFQX1 \a11_reg[4]  ( .D(n1334), .CK(clk), .Q(a11[4]) );
  DFFQX1 \a12_reg[5]  ( .D(n1341), .CK(clk), .Q(a12[5]) );
  DFFQX1 \a12_reg[4]  ( .D(n1342), .CK(clk), .Q(a12[4]) );
  DFFQX1 \a13_reg[5]  ( .D(n1349), .CK(clk), .Q(a13[5]) );
  DFFQX1 \a13_reg[4]  ( .D(n1350), .CK(clk), .Q(a13[4]) );
  DFFX1 \b43_reg[3]  ( .D(n1455), .CK(clk), .Q(b43[3]), .QN(n671) );
  DFFX1 \b43_reg[2]  ( .D(n1456), .CK(clk), .Q(b43[2]), .QN(n672) );
  DFFX1 \b43_reg[1]  ( .D(n1457), .CK(clk), .Q(b43[1]), .QN(n673) );
  DFFX1 \b44_reg[3]  ( .D(n1479), .CK(clk), .Q(b44[3]), .QN(n679) );
  DFFX1 \b44_reg[2]  ( .D(n1480), .CK(clk), .Q(b44[2]), .QN(n680) );
  DFFX1 \b44_reg[1]  ( .D(n1481), .CK(clk), .Q(b44[1]), .QN(n681) );
  DFFX1 \b12_reg[3]  ( .D(n1431), .CK(clk), .Q(b12[3]), .QN(n639) );
  DFFX1 \b12_reg[2]  ( .D(n1432), .CK(clk), .Q(b12[2]), .QN(n640) );
  DFFX1 \b12_reg[1]  ( .D(n1433), .CK(clk), .Q(b12[1]), .QN(n641) );
  DFFX1 \b13_reg[3]  ( .D(n1447), .CK(clk), .Q(b13[3]), .QN(n655) );
  DFFX1 \b13_reg[2]  ( .D(n1448), .CK(clk), .Q(b13[2]), .QN(n656) );
  DFFX1 \b13_reg[1]  ( .D(n1449), .CK(clk), .Q(b13[1]), .QN(n657) );
  DFFX1 \b22_reg[3]  ( .D(n1439), .CK(clk), .Q(b22[3]), .QN(n647) );
  DFFX1 \b22_reg[2]  ( .D(n1440), .CK(clk), .Q(b22[2]), .QN(n648) );
  DFFX1 \b22_reg[1]  ( .D(n1441), .CK(clk), .Q(b22[1]), .QN(n649) );
  DFFX1 \b34_reg[3]  ( .D(n1463), .CK(clk), .Q(b34[3]), .QN(n663) );
  DFFX1 \b34_reg[2]  ( .D(n1464), .CK(clk), .Q(b34[2]), .QN(n664) );
  DFFX1 \b34_reg[1]  ( .D(n1465), .CK(clk), .Q(b34[1]), .QN(n665) );
  DFFX1 \b43_reg[0]  ( .D(n1458), .CK(clk), .Q(b43[0]), .QN(n674) );
  DFFX1 \b44_reg[0]  ( .D(n1482), .CK(clk), .Q(b44[0]), .QN(n682) );
  DFFX1 \b12_reg[0]  ( .D(n1434), .CK(clk), .Q(b12[0]), .QN(n642) );
  DFFX1 \b13_reg[0]  ( .D(n1450), .CK(clk), .Q(b13[0]), .QN(n658) );
  DFFX1 \b22_reg[0]  ( .D(n1442), .CK(clk), .Q(b22[0]), .QN(n650) );
  DFFX1 \b34_reg[0]  ( .D(n1466), .CK(clk), .Q(b34[0]), .QN(n666) );
  DFFQX1 \b41_reg[3]  ( .D(n1423), .CK(clk), .Q(b41[3]) );
  DFFQX1 \b41_reg[2]  ( .D(n1424), .CK(clk), .Q(b41[2]) );
  DFFQX1 \b41_reg[1]  ( .D(n1425), .CK(clk), .Q(b41[1]) );
  DFFQX1 \b11_reg[3]  ( .D(n1399), .CK(clk), .Q(b11[3]) );
  DFFQX1 \b11_reg[2]  ( .D(n1400), .CK(clk), .Q(b11[2]) );
  DFFQX1 \b11_reg[1]  ( .D(n1401), .CK(clk), .Q(b11[1]) );
  DFFQX1 \b21_reg[3]  ( .D(n1407), .CK(clk), .Q(b21[3]) );
  DFFQX1 \b21_reg[2]  ( .D(n1408), .CK(clk), .Q(b21[2]) );
  DFFQX1 \b21_reg[1]  ( .D(n1409), .CK(clk), .Q(b21[1]) );
  DFFQX1 \b31_reg[3]  ( .D(n1415), .CK(clk), .Q(b31[3]) );
  DFFQX1 \b31_reg[2]  ( .D(n1416), .CK(clk), .Q(b31[2]) );
  DFFQX1 \b31_reg[1]  ( .D(n1417), .CK(clk), .Q(b31[1]) );
  DFFQX1 \b42_reg[3]  ( .D(n1877), .CK(clk), .Q(b42[3]) );
  DFFQX1 \b42_reg[2]  ( .D(n1876), .CK(clk), .Q(b42[2]) );
  DFFQX1 \b42_reg[1]  ( .D(n1875), .CK(clk), .Q(b42[1]) );
  DFFQX1 \b14_reg[3]  ( .D(n1885), .CK(clk), .Q(b14[3]) );
  DFFQX1 \b14_reg[2]  ( .D(n1884), .CK(clk), .Q(b14[2]) );
  DFFQX1 \b14_reg[1]  ( .D(n1883), .CK(clk), .Q(b14[1]) );
  DFFQX1 \b23_reg[3]  ( .D(n1893), .CK(clk), .Q(b23[3]) );
  DFFQX1 \b23_reg[2]  ( .D(n1892), .CK(clk), .Q(b23[2]) );
  DFFQX1 \b23_reg[1]  ( .D(n1891), .CK(clk), .Q(b23[1]) );
  DFFQX1 \b24_reg[3]  ( .D(n1861), .CK(clk), .Q(b24[3]) );
  DFFQX1 \b24_reg[2]  ( .D(n1860), .CK(clk), .Q(b24[2]) );
  DFFQX1 \b24_reg[1]  ( .D(n1859), .CK(clk), .Q(b24[1]) );
  DFFQX1 \b32_reg[3]  ( .D(n1901), .CK(clk), .Q(b32[3]) );
  DFFQX1 \b32_reg[2]  ( .D(n1900), .CK(clk), .Q(b32[2]) );
  DFFQX1 \b32_reg[1]  ( .D(n1899), .CK(clk), .Q(b32[1]) );
  DFFQX1 \b33_reg[3]  ( .D(n1869), .CK(clk), .Q(b33[3]) );
  DFFQX1 \b33_reg[2]  ( .D(n1868), .CK(clk), .Q(b33[2]) );
  DFFQX1 \b33_reg[1]  ( .D(n1867), .CK(clk), .Q(b33[1]) );
  DFFQX1 \b41_reg[0]  ( .D(n1426), .CK(clk), .Q(b41[0]) );
  DFFQX1 \b11_reg[0]  ( .D(n1402), .CK(clk), .Q(b11[0]) );
  DFFQX1 \b21_reg[0]  ( .D(n1410), .CK(clk), .Q(b21[0]) );
  DFFQX1 \b31_reg[0]  ( .D(n1418), .CK(clk), .Q(b31[0]) );
  DFFQX1 \a14_reg[3]  ( .D(n1359), .CK(clk), .Q(a14[3]) );
  DFFQX1 \a14_reg[2]  ( .D(n1360), .CK(clk), .Q(a14[2]) );
  DFFQX1 \a14_reg[1]  ( .D(n1361), .CK(clk), .Q(a14[1]) );
  DFFQX1 \a11_reg[3]  ( .D(n1335), .CK(clk), .Q(a11[3]) );
  DFFQX1 \a11_reg[2]  ( .D(n1336), .CK(clk), .Q(a11[2]) );
  DFFQX1 \a11_reg[1]  ( .D(n1337), .CK(clk), .Q(a11[1]) );
  DFFQX1 \a12_reg[3]  ( .D(n1343), .CK(clk), .Q(a12[3]) );
  DFFQX1 \a12_reg[2]  ( .D(n1344), .CK(clk), .Q(a12[2]) );
  DFFQX1 \a12_reg[1]  ( .D(n1345), .CK(clk), .Q(a12[1]) );
  DFFQX1 \a13_reg[3]  ( .D(n1351), .CK(clk), .Q(a13[3]) );
  DFFQX1 \a13_reg[2]  ( .D(n1352), .CK(clk), .Q(a13[2]) );
  DFFQX1 \a13_reg[1]  ( .D(n1353), .CK(clk), .Q(a13[1]) );
  DFFQX1 \b42_reg[0]  ( .D(n1874), .CK(clk), .Q(b42[0]) );
  DFFQX1 \b14_reg[0]  ( .D(n1882), .CK(clk), .Q(b14[0]) );
  DFFQX1 \b23_reg[0]  ( .D(n1890), .CK(clk), .Q(b23[0]) );
  DFFQX1 \b24_reg[0]  ( .D(n1858), .CK(clk), .Q(b24[0]) );
  DFFQX1 \b32_reg[0]  ( .D(n1898), .CK(clk), .Q(b32[0]) );
  DFFQX1 \b33_reg[0]  ( .D(n1866), .CK(clk), .Q(b33[0]) );
  DFFQX1 \a14_reg[0]  ( .D(n1362), .CK(clk), .Q(a14[0]) );
  DFFQX1 \a11_reg[0]  ( .D(n1338), .CK(clk), .Q(a11[0]) );
  DFFQX1 \a12_reg[0]  ( .D(n1346), .CK(clk), .Q(a12[0]) );
  DFFQX1 \a13_reg[0]  ( .D(n1354), .CK(clk), .Q(a13[0]) );
  DFFTRX1 \counter_reg[5]  ( .D(N635), .RN(n1906), .CK(clk), .Q(counter[5]) );
  DFFTRX1 \counter_reg[6]  ( .D(N636), .RN(n1906), .CK(clk), .Q(counter[6]) );
  DFFTRX1 \counter_reg[7]  ( .D(N637), .RN(n1906), .CK(clk), .Q(counter[7]) );
  DFFTRX1 \counter_reg[8]  ( .D(N638), .RN(n1906), .CK(clk), .Q(counter[8]) );
  DFFTRX1 \counter_reg[9]  ( .D(N639), .RN(n1906), .CK(clk), .Q(counter[9]), 
        .QN(n1519) );
  DFFTRX1 \counter_reg[10]  ( .D(N640), .RN(n1906), .CK(clk), .Q(counter[10]), 
        .QN(n1516) );
  DFFTRX1 \counter_reg[2]  ( .D(N632), .RN(n1906), .CK(clk), .Q(counter[2]) );
  DFFTRX1 \counter_reg[3]  ( .D(N633), .RN(n1906), .CK(clk), .Q(counter[3]), 
        .QN(n1515) );
  DFFTRX1 \counter_reg[4]  ( .D(N634), .RN(n1906), .CK(clk), .Q(counter[4]), 
        .QN(n1533) );
  ADDFXL \add_1_root_sub_0_root_sub_359_2/U1_2  ( .A(n[2]), .B(N247), .CI(
        \add_1_root_sub_0_root_sub_359_2/carry[2] ), .CO(
        \add_1_root_sub_0_root_sub_359_2/carry[3] ), .S(N796) );
  ADDFXL \add_1_root_sub_0_root_sub_359_2/U1_1  ( .A(n[1]), .B(N241), .CI(
        n1517), .CO(\add_1_root_sub_0_root_sub_359_2/carry[2] ), .S(N795) );
  ADDFXL \add_1_root_sub_0_root_sub_359_2/U1_3  ( .A(n[3]), .B(k[3]), .CI(
        \add_1_root_sub_0_root_sub_359_2/carry[3] ), .CO(N798), .S(N797) );
  ADDHXL \add_332/U1_1_1  ( .A(N241), .B(N785), .CO(\add_332/carry[2] ), .S(
        N719) );
  ADDHXL \add_332/U1_1_2  ( .A(N247), .B(\add_332/carry[2] ), .CO(
        \add_332/carry[3] ), .S(N720) );
  ADDHXL \add_331/U1_1_1  ( .A(N241), .B(N785), .CO(\add_331/carry[2] ), .S(
        N712) );
  ADDHX1 \add_331/U1_1_3  ( .A(k[3]), .B(\add_331/carry[3] ), .CO(N715), .S(
        N714) );
  DFFQX1 \index_b_reg[5]  ( .D(n1492), .CK(clk), .Q(index_b[5]) );
  DFFQX1 \index_a_reg[5]  ( .D(n1501), .CK(clk), .Q(index_a[5]) );
  DFFQX1 \index_b_reg[6]  ( .D(n1491), .CK(clk), .Q(index_b[6]) );
  DFFQX1 \index_a_reg[6]  ( .D(n1500), .CK(clk), .Q(index_a[6]) );
  DFFTRX1 \counter_reg[1]  ( .D(N631), .RN(n1906), .CK(clk), .Q(counter[1]), 
        .QN(n699) );
  DFFTRX1 \counter_reg[0]  ( .D(N630), .RN(n1906), .CK(clk), .Q(counter[0]), 
        .QN(n700) );
  CMPR32X2 \add_357_2/U1_3  ( .A(k[3]), .B(n[2]), .C(\add_357_2/carry[3] ), 
        .CO(\add_357_2/carry[4] ), .S(N788) );
  DFFXL \temp1_reg[0]  ( .D(n1322), .CK(clk), .QN(n724) );
  DFFXL \temp1_reg[1]  ( .D(n1321), .CK(clk), .QN(n723) );
  DFFXL \temp1_reg[2]  ( .D(n1320), .CK(clk), .QN(n722) );
  DFFXL \temp1_reg[3]  ( .D(n1319), .CK(clk), .QN(n721) );
  DFFXL \temp1_reg[4]  ( .D(n1318), .CK(clk), .QN(n720) );
  DFFXL \temp1_reg[5]  ( .D(n1317), .CK(clk), .QN(n719) );
  DFFXL \temp1_reg[6]  ( .D(n1316), .CK(clk), .QN(n718) );
  DFFXL \temp1_reg[7]  ( .D(n1315), .CK(clk), .QN(n717) );
  DFFXL \temp1_reg[8]  ( .D(n1314), .CK(clk), .QN(n716) );
  DFFXL \temp1_reg[9]  ( .D(n1313), .CK(clk), .QN(n715) );
  DFFXL \temp1_reg[10]  ( .D(n1312), .CK(clk), .QN(n714) );
  DFFXL \temp1_reg[11]  ( .D(n1311), .CK(clk), .QN(n713) );
  DFFXL \temp1_reg[12]  ( .D(n1310), .CK(clk), .QN(n712) );
  DFFXL \temp1_reg[13]  ( .D(n1309), .CK(clk), .QN(n711) );
  DFFXL \temp1_reg[14]  ( .D(n1308), .CK(clk), .QN(n710) );
  DFFXL \temp1_reg[15]  ( .D(n1307), .CK(clk), .QN(n709) );
  EDFFXL \index_out_reg[7]  ( .D(N809), .E(n1680), .CK(clk), .Q(index_out[7])
         );
  EDFFXL \index_out_reg[6]  ( .D(N808), .E(n1680), .CK(clk), .Q(index_out[6])
         );
  DFFXL \temp2_reg[0]  ( .D(n1330), .CK(clk), .QN(n740) );
  DFFXL \temp2_reg[1]  ( .D(n1329), .CK(clk), .QN(n739) );
  DFFXL \temp2_reg[2]  ( .D(n1328), .CK(clk), .QN(n738) );
  DFFXL \temp2_reg[3]  ( .D(n1327), .CK(clk), .QN(n737) );
  DFFXL \temp2_reg[4]  ( .D(n1326), .CK(clk), .QN(n736) );
  DFFXL \temp2_reg[5]  ( .D(n1325), .CK(clk), .QN(n735) );
  DFFXL \temp2_reg[6]  ( .D(n1324), .CK(clk), .QN(n734) );
  DFFXL \temp2_reg[7]  ( .D(n1323), .CK(clk), .QN(n733) );
  DFFQXL \data_in_o_reg[31]  ( .D(n1306), .CK(clk), .Q(data_in_o[31]) );
  DFFQXL \data_in_o_reg[30]  ( .D(n1305), .CK(clk), .Q(data_in_o[30]) );
  DFFQXL \data_in_o_reg[29]  ( .D(n1304), .CK(clk), .Q(data_in_o[29]) );
  DFFQXL \data_in_o_reg[28]  ( .D(n1303), .CK(clk), .Q(data_in_o[28]) );
  DFFQXL \data_in_o_reg[27]  ( .D(n1302), .CK(clk), .Q(data_in_o[27]) );
  DFFQXL \data_in_o_reg[26]  ( .D(n1301), .CK(clk), .Q(data_in_o[26]) );
  DFFQXL \data_in_o_reg[25]  ( .D(n1300), .CK(clk), .Q(data_in_o[25]) );
  DFFQXL \data_in_o_reg[24]  ( .D(n1299), .CK(clk), .Q(data_in_o[24]) );
  DFFQXL \data_in_o_reg[17]  ( .D(n1511), .CK(clk), .Q(data_in_o[17]) );
  DFFQXL \data_in_o_reg[23]  ( .D(n1751), .CK(clk), .Q(data_in_o[23]) );
  DFFQXL \data_in_o_reg[22]  ( .D(n1750), .CK(clk), .Q(data_in_o[22]) );
  DFFQXL \data_in_o_reg[21]  ( .D(n1514), .CK(clk), .Q(data_in_o[21]) );
  DFFQXL \data_in_o_reg[20]  ( .D(n1513), .CK(clk), .Q(data_in_o[20]) );
  DFFQXL \data_in_o_reg[19]  ( .D(n1749), .CK(clk), .Q(data_in_o[19]) );
  DFFQXL \data_in_o_reg[18]  ( .D(n1522), .CK(clk), .Q(data_in_o[18]) );
  DFFQXL \data_in_o_reg[15]  ( .D(n1298), .CK(clk), .Q(data_in_o[15]) );
  DFFQXL \data_in_o_reg[14]  ( .D(n1297), .CK(clk), .Q(data_in_o[14]) );
  DFFQXL \data_in_o_reg[13]  ( .D(n1296), .CK(clk), .Q(data_in_o[13]) );
  DFFQXL \data_in_o_reg[12]  ( .D(n1295), .CK(clk), .Q(data_in_o[12]) );
  DFFQXL \data_in_o_reg[11]  ( .D(n1294), .CK(clk), .Q(data_in_o[11]) );
  DFFQXL \data_in_o_reg[10]  ( .D(n1293), .CK(clk), .Q(data_in_o[10]) );
  DFFQXL \data_in_o_reg[9]  ( .D(n1292), .CK(clk), .Q(data_in_o[9]) );
  DFFQXL \data_in_o_reg[8]  ( .D(n1291), .CK(clk), .Q(data_in_o[8]) );
  DFFQXL \data_in_o_reg[7]  ( .D(n1290), .CK(clk), .Q(data_in_o[7]) );
  DFFQXL \data_in_o_reg[6]  ( .D(n1289), .CK(clk), .Q(data_in_o[6]) );
  DFFQXL \data_in_o_reg[5]  ( .D(n1288), .CK(clk), .Q(data_in_o[5]) );
  DFFQXL \data_in_o_reg[4]  ( .D(n1287), .CK(clk), .Q(data_in_o[4]) );
  DFFQXL \data_in_o_reg[3]  ( .D(n1286), .CK(clk), .Q(data_in_o[3]) );
  DFFQXL \data_in_o_reg[2]  ( .D(n1285), .CK(clk), .Q(data_in_o[2]) );
  DFFQXL \data_in_o_reg[1]  ( .D(n1284), .CK(clk), .Q(data_in_o[1]) );
  DFFQXL \data_in_o_reg[0]  ( .D(n1283), .CK(clk), .Q(data_in_o[0]) );
  ADDFHX4 \add_357/U1_1  ( .A(N241), .B(n[1]), .CI(n1543), .CO(
        \add_357/carry[2] ), .S(N780) );
  DFFQX1 \data_in_o_reg[16]  ( .D(n1512), .CK(clk), .Q(data_in_o[16]) );
  CMPR22X2 \add_331/U1_1_2  ( .A(N247), .B(\add_331/carry[2] ), .CO(
        \add_331/carry[3] ), .S(N713) );
  EDFFXL \l_reg[2]  ( .D(N252), .E(n1907), .CK(clk), .Q(l[2]), .QN(n629) );
  EDFFXL \l_reg[1]  ( .D(N241), .E(n1907), .CK(clk), .Q(l[1]), .QN(n630) );
  EDFFXL \l_reg[0]  ( .D(N785), .E(n1907), .CK(clk), .Q(l[0]), .QN(n631) );
  EDFFXL \matrix_a_reg[8][7]  ( .D(data_out_a[7]), .E(n1560), .CK(clk), .QN(
        n506) );
  EDFFXL \matrix_a_reg[8][6]  ( .D(data_out_a[6]), .E(n1560), .CK(clk), .QN(
        n507) );
  EDFFXL \matrix_a_reg[8][5]  ( .D(data_out_a[5]), .E(n1560), .CK(clk), .QN(
        n508) );
  EDFFXL \matrix_a_reg[8][4]  ( .D(data_out_a[4]), .E(n1560), .CK(clk), .QN(
        n509) );
  EDFFXL \matrix_a_reg[8][3]  ( .D(data_out_a[3]), .E(n1560), .CK(clk), .QN(
        n510) );
  EDFFXL \matrix_a_reg[8][2]  ( .D(data_out_a[2]), .E(n1560), .CK(clk), .QN(
        n511) );
  EDFFXL \matrix_a_reg[8][1]  ( .D(data_out_a[1]), .E(n1560), .CK(clk), .QN(
        n512) );
  EDFFXL \matrix_a_reg[8][0]  ( .D(data_out_a[0]), .E(n1560), .CK(clk), .QN(
        n513) );
  EDFFXL \matrix_a_reg[7][7]  ( .D(data_out_a[7]), .E(n1569), .CK(clk), .QN(
        n474) );
  EDFFXL \matrix_a_reg[7][6]  ( .D(data_out_a[6]), .E(n1569), .CK(clk), .QN(
        n475) );
  EDFFXL \matrix_a_reg[7][5]  ( .D(data_out_a[5]), .E(n1569), .CK(clk), .QN(
        n476) );
  EDFFXL \matrix_a_reg[7][4]  ( .D(data_out_a[4]), .E(n1569), .CK(clk), .QN(
        n477) );
  EDFFXL \matrix_a_reg[7][3]  ( .D(data_out_a[3]), .E(n1569), .CK(clk), .QN(
        n478) );
  EDFFXL \matrix_a_reg[7][2]  ( .D(data_out_a[2]), .E(n1569), .CK(clk), .QN(
        n479) );
  EDFFXL \matrix_a_reg[7][1]  ( .D(data_out_a[1]), .E(n1569), .CK(clk), .QN(
        n480) );
  EDFFXL \matrix_a_reg[7][0]  ( .D(data_out_a[0]), .E(n1569), .CK(clk), .QN(
        n481) );
  EDFFXL \matrix_b_reg[7][7]  ( .D(data_out_b[7]), .E(n1570), .CK(clk), .QN(
        n602) );
  EDFFXL \matrix_b_reg[7][6]  ( .D(data_out_b[6]), .E(n1570), .CK(clk), .QN(
        n603) );
  EDFFXL \matrix_b_reg[7][5]  ( .D(data_out_b[5]), .E(n1570), .CK(clk), .QN(
        n604) );
  EDFFXL \matrix_b_reg[7][4]  ( .D(data_out_b[4]), .E(n1570), .CK(clk), .QN(
        n605) );
  EDFFXL \matrix_b_reg[7][3]  ( .D(data_out_b[3]), .E(n1570), .CK(clk), .QN(
        n606) );
  EDFFXL \matrix_b_reg[7][2]  ( .D(data_out_b[2]), .E(n1570), .CK(clk), .QN(
        n607) );
  EDFFXL \matrix_b_reg[7][1]  ( .D(data_out_b[1]), .E(n1570), .CK(clk), .QN(
        n608) );
  EDFFXL \matrix_b_reg[7][0]  ( .D(data_out_b[0]), .E(n1570), .CK(clk), .QN(
        n609) );
  EDFFXL \matrix_a_reg[8][31]  ( .D(data_out_a[31]), .E(n1560), .CK(clk), .QN(
        n482) );
  EDFFXL \matrix_a_reg[8][30]  ( .D(data_out_a[30]), .E(n1560), .CK(clk), .QN(
        n483) );
  EDFFXL \matrix_a_reg[8][29]  ( .D(data_out_a[29]), .E(n1560), .CK(clk), .QN(
        n484) );
  EDFFXL \matrix_a_reg[8][28]  ( .D(data_out_a[28]), .E(n1560), .CK(clk), .QN(
        n485) );
  EDFFXL \matrix_a_reg[8][27]  ( .D(data_out_a[27]), .E(n1560), .CK(clk), .QN(
        n486) );
  EDFFXL \matrix_a_reg[8][26]  ( .D(data_out_a[26]), .E(n1560), .CK(clk), .QN(
        n487) );
  EDFFXL \matrix_a_reg[8][25]  ( .D(data_out_a[25]), .E(n1560), .CK(clk), .QN(
        n488) );
  EDFFXL \matrix_a_reg[8][24]  ( .D(data_out_a[24]), .E(n1560), .CK(clk), .QN(
        n489) );
  EDFFXL \matrix_a_reg[8][23]  ( .D(data_out_a[23]), .E(n1560), .CK(clk), .QN(
        n490) );
  EDFFXL \matrix_a_reg[8][22]  ( .D(data_out_a[22]), .E(n1560), .CK(clk), .QN(
        n491) );
  EDFFXL \matrix_a_reg[8][21]  ( .D(data_out_a[21]), .E(n1560), .CK(clk), .QN(
        n492) );
  EDFFXL \matrix_a_reg[8][20]  ( .D(data_out_a[20]), .E(n1560), .CK(clk), .QN(
        n493) );
  EDFFXL \matrix_a_reg[8][19]  ( .D(data_out_a[19]), .E(n1560), .CK(clk), .QN(
        n494) );
  EDFFXL \matrix_a_reg[8][18]  ( .D(data_out_a[18]), .E(n1560), .CK(clk), .QN(
        n495) );
  EDFFXL \matrix_a_reg[8][17]  ( .D(data_out_a[17]), .E(n1560), .CK(clk), .QN(
        n496) );
  EDFFXL \matrix_a_reg[8][16]  ( .D(data_out_a[16]), .E(n1560), .CK(clk), .QN(
        n497) );
  EDFFXL \matrix_a_reg[8][15]  ( .D(data_out_a[15]), .E(n1560), .CK(clk), .QN(
        n498) );
  EDFFXL \matrix_a_reg[8][14]  ( .D(data_out_a[14]), .E(n1560), .CK(clk), .QN(
        n499) );
  EDFFXL \matrix_a_reg[8][13]  ( .D(data_out_a[13]), .E(n1560), .CK(clk), .QN(
        n500) );
  EDFFXL \matrix_a_reg[8][12]  ( .D(data_out_a[12]), .E(n1560), .CK(clk), .QN(
        n501) );
  EDFFXL \matrix_a_reg[8][11]  ( .D(data_out_a[11]), .E(n1560), .CK(clk), .QN(
        n502) );
  EDFFXL \matrix_a_reg[8][10]  ( .D(data_out_a[10]), .E(n1560), .CK(clk), .QN(
        n503) );
  EDFFXL \matrix_a_reg[8][9]  ( .D(data_out_a[9]), .E(n1560), .CK(clk), .QN(
        n504) );
  EDFFXL \matrix_a_reg[8][8]  ( .D(data_out_a[8]), .E(n1560), .CK(clk), .QN(
        n505) );
  EDFFXL \matrix_a_reg[7][31]  ( .D(data_out_a[31]), .E(n1569), .CK(clk), .QN(
        n450) );
  EDFFXL \matrix_a_reg[7][30]  ( .D(data_out_a[30]), .E(n1569), .CK(clk), .QN(
        n451) );
  EDFFXL \matrix_a_reg[7][29]  ( .D(data_out_a[29]), .E(n1569), .CK(clk), .QN(
        n452) );
  EDFFXL \matrix_a_reg[7][28]  ( .D(data_out_a[28]), .E(n1569), .CK(clk), .QN(
        n453) );
  EDFFXL \matrix_a_reg[7][27]  ( .D(data_out_a[27]), .E(n1569), .CK(clk), .QN(
        n454) );
  EDFFXL \matrix_a_reg[7][26]  ( .D(data_out_a[26]), .E(n1569), .CK(clk), .QN(
        n455) );
  EDFFXL \matrix_a_reg[7][25]  ( .D(data_out_a[25]), .E(n1569), .CK(clk), .QN(
        n456) );
  EDFFXL \matrix_a_reg[7][24]  ( .D(data_out_a[24]), .E(n1569), .CK(clk), .QN(
        n457) );
  EDFFXL \matrix_b_reg[7][15]  ( .D(data_out_b[15]), .E(n1570), .CK(clk), .QN(
        n594) );
  EDFFXL \matrix_b_reg[7][14]  ( .D(data_out_b[14]), .E(n1570), .CK(clk), .QN(
        n595) );
  EDFFXL \matrix_b_reg[7][13]  ( .D(data_out_b[13]), .E(n1570), .CK(clk), .QN(
        n596) );
  EDFFXL \matrix_b_reg[7][12]  ( .D(data_out_b[12]), .E(n1570), .CK(clk), .QN(
        n597) );
  EDFFXL \matrix_b_reg[7][11]  ( .D(data_out_b[11]), .E(n1570), .CK(clk), .QN(
        n598) );
  EDFFXL \matrix_b_reg[7][10]  ( .D(data_out_b[10]), .E(n1570), .CK(clk), .QN(
        n599) );
  EDFFXL \matrix_b_reg[7][9]  ( .D(data_out_b[9]), .E(n1570), .CK(clk), .QN(
        n600) );
  EDFFXL \matrix_b_reg[7][8]  ( .D(data_out_b[8]), .E(n1570), .CK(clk), .QN(
        n601) );
  EDFFXL \matrix_b_reg[2][7]  ( .D(data_out_b[7]), .E(n1558), .CK(clk), .QN(
        n538) );
  EDFFXL \matrix_b_reg[2][6]  ( .D(data_out_b[6]), .E(n1558), .CK(clk), .QN(
        n539) );
  EDFFXL \matrix_b_reg[2][5]  ( .D(data_out_b[5]), .E(n1558), .CK(clk), .QN(
        n540) );
  EDFFXL \matrix_b_reg[2][4]  ( .D(data_out_b[4]), .E(n1558), .CK(clk), .QN(
        n541) );
  EDFFXL \matrix_b_reg[2][3]  ( .D(data_out_b[3]), .E(n1558), .CK(clk), .QN(
        n542) );
  EDFFXL \matrix_b_reg[2][2]  ( .D(data_out_b[2]), .E(n1558), .CK(clk), .QN(
        n543) );
  EDFFXL \matrix_b_reg[2][1]  ( .D(data_out_b[1]), .E(n1558), .CK(clk), .QN(
        n544) );
  EDFFXL \matrix_b_reg[2][0]  ( .D(data_out_b[0]), .E(n1558), .CK(clk), .QN(
        n545) );
  EDFFXL \matrix_b_reg[5][23]  ( .D(data_out_b[23]), .E(n1563), .CK(clk), .QN(
        n578) );
  EDFFXL \matrix_b_reg[5][22]  ( .D(data_out_b[22]), .E(n1563), .CK(clk), .QN(
        n579) );
  EDFFXL \matrix_b_reg[5][21]  ( .D(data_out_b[21]), .E(n1563), .CK(clk), .QN(
        n580) );
  EDFFXL \matrix_b_reg[5][20]  ( .D(data_out_b[20]), .E(n1563), .CK(clk), .QN(
        n581) );
  EDFFXL \matrix_b_reg[5][19]  ( .D(data_out_b[19]), .E(n1563), .CK(clk), .QN(
        n582) );
  EDFFXL \matrix_b_reg[5][18]  ( .D(data_out_b[18]), .E(n1563), .CK(clk), .QN(
        n583) );
  EDFFXL \matrix_b_reg[5][17]  ( .D(data_out_b[17]), .E(n1563), .CK(clk), .QN(
        n584) );
  EDFFXL \matrix_b_reg[5][16]  ( .D(data_out_b[16]), .E(n1563), .CK(clk), .QN(
        n585) );
  EDFFXL \matrix_b_reg[4][23]  ( .D(data_out_b[23]), .E(n1564), .CK(clk), .QN(
        n562) );
  EDFFXL \matrix_b_reg[4][22]  ( .D(data_out_b[22]), .E(n1564), .CK(clk), .QN(
        n563) );
  EDFFXL \matrix_b_reg[4][21]  ( .D(data_out_b[21]), .E(n1564), .CK(clk), .QN(
        n564) );
  EDFFXL \matrix_b_reg[4][20]  ( .D(data_out_b[20]), .E(n1564), .CK(clk), .QN(
        n565) );
  EDFFXL \matrix_b_reg[4][19]  ( .D(data_out_b[19]), .E(n1564), .CK(clk), .QN(
        n566) );
  EDFFXL \matrix_b_reg[4][18]  ( .D(data_out_b[18]), .E(n1564), .CK(clk), .QN(
        n567) );
  EDFFXL \matrix_b_reg[4][17]  ( .D(data_out_b[17]), .E(n1564), .CK(clk), .QN(
        n568) );
  EDFFXL \matrix_b_reg[4][16]  ( .D(data_out_b[16]), .E(n1564), .CK(clk), .QN(
        n569) );
  EDFFXL \matrix_b_reg[4][15]  ( .D(data_out_b[15]), .E(n1564), .CK(clk), .QN(
        n570) );
  EDFFXL \matrix_b_reg[4][14]  ( .D(data_out_b[14]), .E(n1564), .CK(clk), .QN(
        n571) );
  EDFFXL \matrix_b_reg[4][13]  ( .D(data_out_b[13]), .E(n1564), .CK(clk), .QN(
        n572) );
  EDFFXL \matrix_b_reg[4][12]  ( .D(data_out_b[12]), .E(n1564), .CK(clk), .QN(
        n573) );
  EDFFXL \matrix_b_reg[4][11]  ( .D(data_out_b[11]), .E(n1564), .CK(clk), .QN(
        n574) );
  EDFFXL \matrix_b_reg[4][10]  ( .D(data_out_b[10]), .E(n1564), .CK(clk), .QN(
        n575) );
  EDFFXL \matrix_b_reg[4][9]  ( .D(data_out_b[9]), .E(n1564), .CK(clk), .QN(
        n576) );
  EDFFXL \matrix_b_reg[4][8]  ( .D(data_out_b[8]), .E(n1564), .CK(clk), .QN(
        n577) );
  EDFFXL \matrix_b_reg[2][31]  ( .D(data_out_b[31]), .E(n1558), .CK(clk), .QN(
        n530) );
  EDFFXL \matrix_b_reg[2][30]  ( .D(data_out_b[30]), .E(n1558), .CK(clk), .QN(
        n531) );
  EDFFXL \matrix_b_reg[2][29]  ( .D(data_out_b[29]), .E(n1558), .CK(clk), .QN(
        n532) );
  EDFFXL \matrix_b_reg[2][28]  ( .D(data_out_b[28]), .E(n1558), .CK(clk), .QN(
        n533) );
  EDFFXL \matrix_b_reg[2][27]  ( .D(data_out_b[27]), .E(n1558), .CK(clk), .QN(
        n534) );
  EDFFXL \matrix_b_reg[2][26]  ( .D(data_out_b[26]), .E(n1558), .CK(clk), .QN(
        n535) );
  EDFFXL \matrix_b_reg[2][25]  ( .D(data_out_b[25]), .E(n1558), .CK(clk), .QN(
        n536) );
  EDFFXL \matrix_b_reg[2][24]  ( .D(data_out_b[24]), .E(n1558), .CK(clk), .QN(
        n537) );
  EDFFXL \matrix_b_reg[1][31]  ( .D(data_out_b[31]), .E(n1567), .CK(clk), .QN(
        n514) );
  EDFFXL \matrix_b_reg[1][30]  ( .D(data_out_b[30]), .E(n1567), .CK(clk), .QN(
        n515) );
  EDFFXL \matrix_b_reg[1][29]  ( .D(data_out_b[29]), .E(n1567), .CK(clk), .QN(
        n516) );
  EDFFXL \matrix_b_reg[1][28]  ( .D(data_out_b[28]), .E(n1567), .CK(clk), .QN(
        n517) );
  EDFFXL \matrix_b_reg[1][27]  ( .D(data_out_b[27]), .E(n1567), .CK(clk), .QN(
        n518) );
  EDFFXL \matrix_b_reg[1][26]  ( .D(data_out_b[26]), .E(n1567), .CK(clk), .QN(
        n519) );
  EDFFXL \matrix_b_reg[1][25]  ( .D(data_out_b[25]), .E(n1567), .CK(clk), .QN(
        n520) );
  EDFFXL \matrix_b_reg[1][24]  ( .D(data_out_b[24]), .E(n1567), .CK(clk), .QN(
        n521) );
  EDFFXL \matrix_b_reg[1][23]  ( .D(data_out_b[23]), .E(n1567), .CK(clk), .QN(
        n522) );
  EDFFXL \matrix_b_reg[1][22]  ( .D(data_out_b[22]), .E(n1567), .CK(clk), .QN(
        n523) );
  EDFFXL \matrix_b_reg[1][21]  ( .D(data_out_b[21]), .E(n1567), .CK(clk), .QN(
        n524) );
  EDFFXL \matrix_b_reg[1][20]  ( .D(data_out_b[20]), .E(n1567), .CK(clk), .QN(
        n525) );
  EDFFXL \matrix_b_reg[1][19]  ( .D(data_out_b[19]), .E(n1567), .CK(clk), .QN(
        n526) );
  EDFFXL \matrix_b_reg[1][18]  ( .D(data_out_b[18]), .E(n1567), .CK(clk), .QN(
        n527) );
  EDFFXL \matrix_b_reg[1][17]  ( .D(data_out_b[17]), .E(n1567), .CK(clk), .QN(
        n528) );
  EDFFXL \matrix_b_reg[1][16]  ( .D(data_out_b[16]), .E(n1567), .CK(clk), .QN(
        n529) );
  EDFFXL \matrix_b_reg[8][19]  ( .D(data_out_b[19]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][19] ) );
  EDFFXL \matrix_b_reg[8][18]  ( .D(data_out_b[18]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][18] ) );
  EDFFXL \matrix_b_reg[8][17]  ( .D(data_out_b[17]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][17] ) );
  EDFFXL \matrix_b_reg[8][16]  ( .D(data_out_b[16]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][16] ) );
  EDFFXL \matrix_b_reg[7][31]  ( .D(data_out_b[31]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][31] ) );
  EDFFXL \matrix_b_reg[7][30]  ( .D(data_out_b[30]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][30] ) );
  EDFFXL \matrix_b_reg[7][29]  ( .D(data_out_b[29]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][29] ) );
  EDFFXL \matrix_b_reg[7][28]  ( .D(data_out_b[28]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][28] ) );
  EDFFXL \matrix_b_reg[7][27]  ( .D(data_out_b[27]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][27] ) );
  EDFFXL \matrix_b_reg[7][26]  ( .D(data_out_b[26]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][26] ) );
  EDFFXL \matrix_b_reg[7][25]  ( .D(data_out_b[25]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][25] ) );
  EDFFXL \matrix_b_reg[7][24]  ( .D(data_out_b[24]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][24] ) );
  EDFFXL \matrix_b_reg[7][19]  ( .D(data_out_b[19]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][19] ) );
  EDFFXL \matrix_b_reg[7][18]  ( .D(data_out_b[18]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][18] ) );
  EDFFXL \matrix_b_reg[7][17]  ( .D(data_out_b[17]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][17] ) );
  EDFFXL \matrix_b_reg[7][16]  ( .D(data_out_b[16]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][16] ) );
  EDFFXL \matrix_b_reg[0][19]  ( .D(data_out_b[19]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][19] ) );
  EDFFXL \matrix_b_reg[0][18]  ( .D(data_out_b[18]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][18] ) );
  EDFFXL \matrix_b_reg[0][17]  ( .D(data_out_b[17]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][17] ) );
  EDFFXL \matrix_b_reg[0][16]  ( .D(data_out_b[16]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][16] ) );
  EDFFXL \matrix_b_reg[6][19]  ( .D(data_out_b[19]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][19] ) );
  EDFFXL \matrix_b_reg[6][18]  ( .D(data_out_b[18]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][18] ) );
  EDFFXL \matrix_b_reg[6][17]  ( .D(data_out_b[17]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][17] ) );
  EDFFXL \matrix_b_reg[6][16]  ( .D(data_out_b[16]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][16] ) );
  EDFFXL \matrix_b_reg[2][19]  ( .D(data_out_b[19]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][19] ) );
  EDFFXL \matrix_b_reg[2][18]  ( .D(data_out_b[18]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][18] ) );
  EDFFXL \matrix_b_reg[2][17]  ( .D(data_out_b[17]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][17] ) );
  EDFFXL \matrix_b_reg[2][16]  ( .D(data_out_b[16]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][16] ) );
  EDFFXL \matrix_b_reg[3][16]  ( .D(data_out_b[16]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][16] ) );
  EDFFXL \matrix_b_reg[3][19]  ( .D(data_out_b[19]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][19] ) );
  EDFFXL \matrix_b_reg[3][18]  ( .D(data_out_b[18]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][18] ) );
  EDFFXL \matrix_b_reg[3][17]  ( .D(data_out_b[17]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][17] ) );
  EDFFX1 \matrix_a_reg[0][31]  ( .D(data_out_a[31]), .E(n1547), .CK(clk), .QN(
        n226) );
  EDFFX1 \matrix_a_reg[5][31]  ( .D(data_out_a[31]), .E(n1565), .CK(clk), .QN(
        n386) );
  EDFFX1 \matrix_a_reg[4][31]  ( .D(data_out_a[31]), .E(n1566), .CK(clk), .QN(
        n354) );
  EDFFX1 \matrix_a_reg[2][31]  ( .D(data_out_a[31]), .E(n1559), .CK(clk), .QN(
        n290) );
  EDFFX1 \matrix_a_reg[1][31]  ( .D(data_out_a[31]), .E(n1568), .CK(clk), .QN(
        n258) );
  EDFFX1 \matrix_a_reg[0][30]  ( .D(data_out_a[30]), .E(n1547), .CK(clk), .QN(
        n227) );
  EDFFX1 \matrix_a_reg[5][30]  ( .D(data_out_a[30]), .E(n1565), .CK(clk), .QN(
        n387) );
  EDFFX1 \matrix_a_reg[4][30]  ( .D(data_out_a[30]), .E(n1566), .CK(clk), .QN(
        n355) );
  EDFFX1 \matrix_a_reg[2][30]  ( .D(data_out_a[30]), .E(n1559), .CK(clk), .QN(
        n291) );
  EDFFX1 \matrix_a_reg[1][30]  ( .D(data_out_a[30]), .E(n1568), .CK(clk), .QN(
        n259) );
  EDFFX1 \matrix_a_reg[0][29]  ( .D(data_out_a[29]), .E(n1547), .CK(clk), .QN(
        n228) );
  EDFFX1 \matrix_a_reg[5][29]  ( .D(data_out_a[29]), .E(n1565), .CK(clk), .QN(
        n388) );
  EDFFX1 \matrix_a_reg[4][29]  ( .D(data_out_a[29]), .E(n1566), .CK(clk), .QN(
        n356) );
  EDFFX1 \matrix_a_reg[2][29]  ( .D(data_out_a[29]), .E(n1559), .CK(clk), .QN(
        n292) );
  EDFFX1 \matrix_a_reg[1][29]  ( .D(data_out_a[29]), .E(n1568), .CK(clk), .QN(
        n260) );
  EDFFX1 \matrix_a_reg[0][28]  ( .D(data_out_a[28]), .E(n1547), .CK(clk), .QN(
        n229) );
  EDFFX1 \matrix_a_reg[5][28]  ( .D(data_out_a[28]), .E(n1565), .CK(clk), .QN(
        n389) );
  EDFFX1 \matrix_a_reg[4][28]  ( .D(data_out_a[28]), .E(n1566), .CK(clk), .QN(
        n357) );
  EDFFX1 \matrix_a_reg[2][28]  ( .D(data_out_a[28]), .E(n1559), .CK(clk), .QN(
        n293) );
  EDFFX1 \matrix_a_reg[1][28]  ( .D(data_out_a[28]), .E(n1568), .CK(clk), .QN(
        n261) );
  EDFFX1 \matrix_a_reg[0][27]  ( .D(data_out_a[27]), .E(n1547), .CK(clk), .QN(
        n230) );
  EDFFX1 \matrix_a_reg[5][27]  ( .D(data_out_a[27]), .E(n1565), .CK(clk), .QN(
        n390) );
  EDFFX1 \matrix_a_reg[4][27]  ( .D(data_out_a[27]), .E(n1566), .CK(clk), .QN(
        n358) );
  EDFFX1 \matrix_a_reg[2][27]  ( .D(data_out_a[27]), .E(n1559), .CK(clk), .QN(
        n294) );
  EDFFX1 \matrix_a_reg[1][27]  ( .D(data_out_a[27]), .E(n1568), .CK(clk), .QN(
        n262) );
  EDFFX1 \matrix_a_reg[0][26]  ( .D(data_out_a[26]), .E(n1547), .CK(clk), .QN(
        n231) );
  EDFFX1 \matrix_a_reg[5][26]  ( .D(data_out_a[26]), .E(n1565), .CK(clk), .QN(
        n391) );
  EDFFX1 \matrix_a_reg[4][26]  ( .D(data_out_a[26]), .E(n1566), .CK(clk), .QN(
        n359) );
  EDFFX1 \matrix_a_reg[2][26]  ( .D(data_out_a[26]), .E(n1559), .CK(clk), .QN(
        n295) );
  EDFFX1 \matrix_a_reg[1][26]  ( .D(data_out_a[26]), .E(n1568), .CK(clk), .QN(
        n263) );
  EDFFX1 \matrix_a_reg[0][25]  ( .D(data_out_a[25]), .E(n1547), .CK(clk), .QN(
        n232) );
  EDFFX1 \matrix_a_reg[5][25]  ( .D(data_out_a[25]), .E(n1565), .CK(clk), .QN(
        n392) );
  EDFFX1 \matrix_a_reg[4][25]  ( .D(data_out_a[25]), .E(n1566), .CK(clk), .QN(
        n360) );
  EDFFX1 \matrix_a_reg[2][25]  ( .D(data_out_a[25]), .E(n1559), .CK(clk), .QN(
        n296) );
  EDFFX1 \matrix_a_reg[1][25]  ( .D(data_out_a[25]), .E(n1568), .CK(clk), .QN(
        n264) );
  EDFFX1 \matrix_a_reg[0][24]  ( .D(data_out_a[24]), .E(n1547), .CK(clk), .QN(
        n233) );
  EDFFX1 \matrix_a_reg[5][24]  ( .D(data_out_a[24]), .E(n1565), .CK(clk), .QN(
        n393) );
  EDFFX1 \matrix_a_reg[4][24]  ( .D(data_out_a[24]), .E(n1566), .CK(clk), .QN(
        n361) );
  EDFFX1 \matrix_a_reg[2][24]  ( .D(data_out_a[24]), .E(n1559), .CK(clk), .QN(
        n297) );
  EDFFX1 \matrix_a_reg[1][24]  ( .D(data_out_a[24]), .E(n1568), .CK(clk), .QN(
        n265) );
  EDFFX1 \matrix_a_reg[0][7]  ( .D(data_out_a[7]), .E(n1547), .CK(clk), .QN(
        n250) );
  EDFFX1 \matrix_a_reg[5][7]  ( .D(data_out_a[7]), .E(n1565), .CK(clk), .QN(
        n410) );
  EDFFX1 \matrix_a_reg[4][7]  ( .D(data_out_a[7]), .E(n1566), .CK(clk), .QN(
        n378) );
  EDFFX1 \matrix_a_reg[2][7]  ( .D(data_out_a[7]), .E(n1559), .CK(clk), .QN(
        n314) );
  EDFFX1 \matrix_a_reg[1][7]  ( .D(data_out_a[7]), .E(n1568), .CK(clk), .QN(
        n282) );
  EDFFX1 \matrix_a_reg[0][6]  ( .D(data_out_a[6]), .E(n1547), .CK(clk), .QN(
        n251) );
  EDFFX1 \matrix_a_reg[5][6]  ( .D(data_out_a[6]), .E(n1565), .CK(clk), .QN(
        n411) );
  EDFFX1 \matrix_a_reg[4][6]  ( .D(data_out_a[6]), .E(n1566), .CK(clk), .QN(
        n379) );
  EDFFX1 \matrix_a_reg[2][6]  ( .D(data_out_a[6]), .E(n1559), .CK(clk), .QN(
        n315) );
  EDFFX1 \matrix_a_reg[1][6]  ( .D(data_out_a[6]), .E(n1568), .CK(clk), .QN(
        n283) );
  EDFFX1 \matrix_a_reg[0][5]  ( .D(data_out_a[5]), .E(n1547), .CK(clk), .QN(
        n252) );
  EDFFX1 \matrix_a_reg[5][5]  ( .D(data_out_a[5]), .E(n1565), .CK(clk), .QN(
        n412) );
  EDFFX1 \matrix_a_reg[4][5]  ( .D(data_out_a[5]), .E(n1566), .CK(clk), .QN(
        n380) );
  EDFFX1 \matrix_a_reg[2][5]  ( .D(data_out_a[5]), .E(n1559), .CK(clk), .QN(
        n316) );
  EDFFX1 \matrix_a_reg[1][5]  ( .D(data_out_a[5]), .E(n1568), .CK(clk), .QN(
        n284) );
  EDFFX1 \matrix_a_reg[0][4]  ( .D(data_out_a[4]), .E(n1547), .CK(clk), .QN(
        n253) );
  EDFFX1 \matrix_a_reg[5][4]  ( .D(data_out_a[4]), .E(n1565), .CK(clk), .QN(
        n413) );
  EDFFX1 \matrix_a_reg[4][4]  ( .D(data_out_a[4]), .E(n1566), .CK(clk), .QN(
        n381) );
  EDFFX1 \matrix_a_reg[2][4]  ( .D(data_out_a[4]), .E(n1559), .CK(clk), .QN(
        n317) );
  EDFFX1 \matrix_a_reg[1][4]  ( .D(data_out_a[4]), .E(n1568), .CK(clk), .QN(
        n285) );
  EDFFX1 \matrix_a_reg[0][3]  ( .D(data_out_a[3]), .E(n1547), .CK(clk), .QN(
        n254) );
  EDFFX1 \matrix_a_reg[5][3]  ( .D(data_out_a[3]), .E(n1565), .CK(clk), .QN(
        n414) );
  EDFFX1 \matrix_a_reg[4][3]  ( .D(data_out_a[3]), .E(n1566), .CK(clk), .QN(
        n382) );
  EDFFX1 \matrix_a_reg[2][3]  ( .D(data_out_a[3]), .E(n1559), .CK(clk), .QN(
        n318) );
  EDFFX1 \matrix_a_reg[1][3]  ( .D(data_out_a[3]), .E(n1568), .CK(clk), .QN(
        n286) );
  EDFFX1 \matrix_a_reg[0][2]  ( .D(data_out_a[2]), .E(n1547), .CK(clk), .QN(
        n255) );
  EDFFX1 \matrix_a_reg[5][2]  ( .D(data_out_a[2]), .E(n1565), .CK(clk), .QN(
        n415) );
  EDFFX1 \matrix_a_reg[4][2]  ( .D(data_out_a[2]), .E(n1566), .CK(clk), .QN(
        n383) );
  EDFFX1 \matrix_a_reg[2][2]  ( .D(data_out_a[2]), .E(n1559), .CK(clk), .QN(
        n319) );
  EDFFX1 \matrix_a_reg[1][2]  ( .D(data_out_a[2]), .E(n1568), .CK(clk), .QN(
        n287) );
  EDFFX1 \matrix_a_reg[0][1]  ( .D(data_out_a[1]), .E(n1547), .CK(clk), .QN(
        n256) );
  EDFFX1 \matrix_a_reg[5][1]  ( .D(data_out_a[1]), .E(n1565), .CK(clk), .QN(
        n416) );
  EDFFX1 \matrix_a_reg[4][1]  ( .D(data_out_a[1]), .E(n1566), .CK(clk), .QN(
        n384) );
  EDFFX1 \matrix_a_reg[2][1]  ( .D(data_out_a[1]), .E(n1559), .CK(clk), .QN(
        n320) );
  EDFFX1 \matrix_a_reg[1][1]  ( .D(data_out_a[1]), .E(n1568), .CK(clk), .QN(
        n288) );
  EDFFX1 \matrix_a_reg[0][0]  ( .D(data_out_a[0]), .E(n1547), .CK(clk), .QN(
        n257) );
  EDFFX1 \matrix_a_reg[5][0]  ( .D(data_out_a[0]), .E(n1565), .CK(clk), .QN(
        n417) );
  EDFFX1 \matrix_a_reg[4][0]  ( .D(data_out_a[0]), .E(n1566), .CK(clk), .QN(
        n385) );
  EDFFX1 \matrix_a_reg[2][0]  ( .D(data_out_a[0]), .E(n1559), .CK(clk), .QN(
        n321) );
  EDFFX1 \matrix_a_reg[1][0]  ( .D(data_out_a[0]), .E(n1568), .CK(clk), .QN(
        n289) );
  EDFFX1 \matrix_a_reg[7][23]  ( .D(data_out_a[23]), .E(n1569), .CK(clk), .QN(
        n458) );
  EDFFX1 \matrix_a_reg[0][23]  ( .D(data_out_a[23]), .E(n1547), .CK(clk), .QN(
        n234) );
  EDFFX1 \matrix_a_reg[5][23]  ( .D(data_out_a[23]), .E(n1565), .CK(clk), .QN(
        n394) );
  EDFFX1 \matrix_a_reg[4][23]  ( .D(data_out_a[23]), .E(n1566), .CK(clk), .QN(
        n362) );
  EDFFX1 \matrix_a_reg[2][23]  ( .D(data_out_a[23]), .E(n1559), .CK(clk), .QN(
        n298) );
  EDFFX1 \matrix_a_reg[7][22]  ( .D(data_out_a[22]), .E(n1569), .CK(clk), .QN(
        n459) );
  EDFFX1 \matrix_a_reg[0][22]  ( .D(data_out_a[22]), .E(n1547), .CK(clk), .QN(
        n235) );
  EDFFX1 \matrix_a_reg[5][22]  ( .D(data_out_a[22]), .E(n1565), .CK(clk), .QN(
        n395) );
  EDFFX1 \matrix_a_reg[4][22]  ( .D(data_out_a[22]), .E(n1566), .CK(clk), .QN(
        n363) );
  EDFFX1 \matrix_a_reg[2][22]  ( .D(data_out_a[22]), .E(n1559), .CK(clk), .QN(
        n299) );
  EDFFX1 \matrix_a_reg[7][21]  ( .D(data_out_a[21]), .E(n1569), .CK(clk), .QN(
        n460) );
  EDFFX1 \matrix_a_reg[0][21]  ( .D(data_out_a[21]), .E(n1547), .CK(clk), .QN(
        n236) );
  EDFFX1 \matrix_a_reg[5][21]  ( .D(data_out_a[21]), .E(n1565), .CK(clk), .QN(
        n396) );
  EDFFX1 \matrix_a_reg[4][21]  ( .D(data_out_a[21]), .E(n1566), .CK(clk), .QN(
        n364) );
  EDFFX1 \matrix_a_reg[2][21]  ( .D(data_out_a[21]), .E(n1559), .CK(clk), .QN(
        n300) );
  EDFFX1 \matrix_a_reg[7][20]  ( .D(data_out_a[20]), .E(n1569), .CK(clk), .QN(
        n461) );
  EDFFX1 \matrix_a_reg[0][20]  ( .D(data_out_a[20]), .E(n1547), .CK(clk), .QN(
        n237) );
  EDFFX1 \matrix_a_reg[5][20]  ( .D(data_out_a[20]), .E(n1565), .CK(clk), .QN(
        n397) );
  EDFFX1 \matrix_a_reg[4][20]  ( .D(data_out_a[20]), .E(n1566), .CK(clk), .QN(
        n365) );
  EDFFX1 \matrix_a_reg[2][20]  ( .D(data_out_a[20]), .E(n1559), .CK(clk), .QN(
        n301) );
  EDFFX1 \matrix_a_reg[7][19]  ( .D(data_out_a[19]), .E(n1569), .CK(clk), .QN(
        n462) );
  EDFFX1 \matrix_a_reg[0][19]  ( .D(data_out_a[19]), .E(n1547), .CK(clk), .QN(
        n238) );
  EDFFX1 \matrix_a_reg[5][19]  ( .D(data_out_a[19]), .E(n1565), .CK(clk), .QN(
        n398) );
  EDFFX1 \matrix_a_reg[4][19]  ( .D(data_out_a[19]), .E(n1566), .CK(clk), .QN(
        n366) );
  EDFFX1 \matrix_a_reg[2][19]  ( .D(data_out_a[19]), .E(n1559), .CK(clk), .QN(
        n302) );
  EDFFX1 \matrix_a_reg[7][18]  ( .D(data_out_a[18]), .E(n1569), .CK(clk), .QN(
        n463) );
  EDFFX1 \matrix_a_reg[0][18]  ( .D(data_out_a[18]), .E(n1547), .CK(clk), .QN(
        n239) );
  EDFFX1 \matrix_a_reg[5][18]  ( .D(data_out_a[18]), .E(n1565), .CK(clk), .QN(
        n399) );
  EDFFX1 \matrix_a_reg[4][18]  ( .D(data_out_a[18]), .E(n1566), .CK(clk), .QN(
        n367) );
  EDFFX1 \matrix_a_reg[2][18]  ( .D(data_out_a[18]), .E(n1559), .CK(clk), .QN(
        n303) );
  EDFFX1 \matrix_a_reg[7][17]  ( .D(data_out_a[17]), .E(n1569), .CK(clk), .QN(
        n464) );
  EDFFX1 \matrix_a_reg[0][17]  ( .D(data_out_a[17]), .E(n1547), .CK(clk), .QN(
        n240) );
  EDFFX1 \matrix_a_reg[5][17]  ( .D(data_out_a[17]), .E(n1565), .CK(clk), .QN(
        n400) );
  EDFFX1 \matrix_a_reg[4][17]  ( .D(data_out_a[17]), .E(n1566), .CK(clk), .QN(
        n368) );
  EDFFX1 \matrix_a_reg[2][17]  ( .D(data_out_a[17]), .E(n1559), .CK(clk), .QN(
        n304) );
  EDFFX1 \matrix_a_reg[7][16]  ( .D(data_out_a[16]), .E(n1569), .CK(clk), .QN(
        n465) );
  EDFFX1 \matrix_a_reg[0][16]  ( .D(data_out_a[16]), .E(n1547), .CK(clk), .QN(
        n241) );
  EDFFX1 \matrix_a_reg[5][16]  ( .D(data_out_a[16]), .E(n1565), .CK(clk), .QN(
        n401) );
  EDFFX1 \matrix_a_reg[4][16]  ( .D(data_out_a[16]), .E(n1566), .CK(clk), .QN(
        n369) );
  EDFFX1 \matrix_a_reg[2][16]  ( .D(data_out_a[16]), .E(n1559), .CK(clk), .QN(
        n305) );
  EDFFX1 \matrix_a_reg[7][15]  ( .D(data_out_a[15]), .E(n1569), .CK(clk), .QN(
        n466) );
  EDFFX1 \matrix_a_reg[0][15]  ( .D(data_out_a[15]), .E(n1547), .CK(clk), .QN(
        n242) );
  EDFFX1 \matrix_a_reg[5][15]  ( .D(data_out_a[15]), .E(n1565), .CK(clk), .QN(
        n402) );
  EDFFX1 \matrix_a_reg[4][15]  ( .D(data_out_a[15]), .E(n1566), .CK(clk), .QN(
        n370) );
  EDFFX1 \matrix_a_reg[2][15]  ( .D(data_out_a[15]), .E(n1559), .CK(clk), .QN(
        n306) );
  EDFFX1 \matrix_a_reg[7][14]  ( .D(data_out_a[14]), .E(n1569), .CK(clk), .QN(
        n467) );
  EDFFX1 \matrix_a_reg[0][14]  ( .D(data_out_a[14]), .E(n1547), .CK(clk), .QN(
        n243) );
  EDFFX1 \matrix_a_reg[5][14]  ( .D(data_out_a[14]), .E(n1565), .CK(clk), .QN(
        n403) );
  EDFFX1 \matrix_a_reg[4][14]  ( .D(data_out_a[14]), .E(n1566), .CK(clk), .QN(
        n371) );
  EDFFX1 \matrix_a_reg[2][14]  ( .D(data_out_a[14]), .E(n1559), .CK(clk), .QN(
        n307) );
  EDFFX1 \matrix_a_reg[7][13]  ( .D(data_out_a[13]), .E(n1569), .CK(clk), .QN(
        n468) );
  EDFFX1 \matrix_a_reg[0][13]  ( .D(data_out_a[13]), .E(n1547), .CK(clk), .QN(
        n244) );
  EDFFX1 \matrix_a_reg[5][13]  ( .D(data_out_a[13]), .E(n1565), .CK(clk), .QN(
        n404) );
  EDFFX1 \matrix_a_reg[4][13]  ( .D(data_out_a[13]), .E(n1566), .CK(clk), .QN(
        n372) );
  EDFFX1 \matrix_a_reg[2][13]  ( .D(data_out_a[13]), .E(n1559), .CK(clk), .QN(
        n308) );
  EDFFX1 \matrix_a_reg[7][12]  ( .D(data_out_a[12]), .E(n1569), .CK(clk), .QN(
        n469) );
  EDFFX1 \matrix_a_reg[0][12]  ( .D(data_out_a[12]), .E(n1547), .CK(clk), .QN(
        n245) );
  EDFFX1 \matrix_a_reg[5][12]  ( .D(data_out_a[12]), .E(n1565), .CK(clk), .QN(
        n405) );
  EDFFX1 \matrix_a_reg[4][12]  ( .D(data_out_a[12]), .E(n1566), .CK(clk), .QN(
        n373) );
  EDFFX1 \matrix_a_reg[2][12]  ( .D(data_out_a[12]), .E(n1559), .CK(clk), .QN(
        n309) );
  EDFFX1 \matrix_a_reg[7][11]  ( .D(data_out_a[11]), .E(n1569), .CK(clk), .QN(
        n470) );
  EDFFX1 \matrix_a_reg[0][11]  ( .D(data_out_a[11]), .E(n1547), .CK(clk), .QN(
        n246) );
  EDFFX1 \matrix_a_reg[5][11]  ( .D(data_out_a[11]), .E(n1565), .CK(clk), .QN(
        n406) );
  EDFFX1 \matrix_a_reg[4][11]  ( .D(data_out_a[11]), .E(n1566), .CK(clk), .QN(
        n374) );
  EDFFX1 \matrix_a_reg[2][11]  ( .D(data_out_a[11]), .E(n1559), .CK(clk), .QN(
        n310) );
  EDFFX1 \matrix_a_reg[7][10]  ( .D(data_out_a[10]), .E(n1569), .CK(clk), .QN(
        n471) );
  EDFFX1 \matrix_a_reg[0][10]  ( .D(data_out_a[10]), .E(n1547), .CK(clk), .QN(
        n247) );
  EDFFX1 \matrix_a_reg[5][10]  ( .D(data_out_a[10]), .E(n1565), .CK(clk), .QN(
        n407) );
  EDFFX1 \matrix_a_reg[4][10]  ( .D(data_out_a[10]), .E(n1566), .CK(clk), .QN(
        n375) );
  EDFFX1 \matrix_a_reg[2][10]  ( .D(data_out_a[10]), .E(n1559), .CK(clk), .QN(
        n311) );
  EDFFX1 \matrix_a_reg[7][9]  ( .D(data_out_a[9]), .E(n1569), .CK(clk), .QN(
        n472) );
  EDFFX1 \matrix_a_reg[0][9]  ( .D(data_out_a[9]), .E(n1547), .CK(clk), .QN(
        n248) );
  EDFFX1 \matrix_a_reg[5][9]  ( .D(data_out_a[9]), .E(n1565), .CK(clk), .QN(
        n408) );
  EDFFX1 \matrix_a_reg[4][9]  ( .D(data_out_a[9]), .E(n1566), .CK(clk), .QN(
        n376) );
  EDFFX1 \matrix_a_reg[2][9]  ( .D(data_out_a[9]), .E(n1559), .CK(clk), .QN(
        n312) );
  EDFFX1 \matrix_a_reg[7][8]  ( .D(data_out_a[8]), .E(n1569), .CK(clk), .QN(
        n473) );
  EDFFX1 \matrix_a_reg[0][8]  ( .D(data_out_a[8]), .E(n1547), .CK(clk), .QN(
        n249) );
  EDFFX1 \matrix_a_reg[5][8]  ( .D(data_out_a[8]), .E(n1565), .CK(clk), .QN(
        n409) );
  EDFFX1 \matrix_a_reg[4][8]  ( .D(data_out_a[8]), .E(n1566), .CK(clk), .QN(
        n377) );
  EDFFX1 \matrix_a_reg[2][8]  ( .D(data_out_a[8]), .E(n1559), .CK(clk), .QN(
        n313) );
  EDFFX1 \matrix_b_reg[0][31]  ( .D(data_out_b[31]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][31] ) );
  EDFFX1 \matrix_b_reg[8][31]  ( .D(data_out_b[31]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][31] ) );
  EDFFX1 \matrix_b_reg[6][31]  ( .D(data_out_b[31]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][31] ) );
  EDFFX1 \matrix_b_reg[5][31]  ( .D(data_out_b[31]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][31] ) );
  EDFFX1 \matrix_b_reg[4][31]  ( .D(data_out_b[31]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][31] ) );
  EDFFX1 \matrix_b_reg[3][31]  ( .D(data_out_b[31]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][31] ) );
  EDFFX1 \matrix_b_reg[0][30]  ( .D(data_out_b[30]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][30] ) );
  EDFFX1 \matrix_b_reg[8][30]  ( .D(data_out_b[30]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][30] ) );
  EDFFX1 \matrix_b_reg[6][30]  ( .D(data_out_b[30]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][30] ) );
  EDFFX1 \matrix_b_reg[5][30]  ( .D(data_out_b[30]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][30] ) );
  EDFFX1 \matrix_b_reg[4][30]  ( .D(data_out_b[30]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][30] ) );
  EDFFX1 \matrix_b_reg[3][30]  ( .D(data_out_b[30]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][30] ) );
  EDFFX1 \matrix_b_reg[0][29]  ( .D(data_out_b[29]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][29] ) );
  EDFFX1 \matrix_b_reg[8][29]  ( .D(data_out_b[29]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][29] ) );
  EDFFX1 \matrix_b_reg[6][29]  ( .D(data_out_b[29]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][29] ) );
  EDFFX1 \matrix_b_reg[5][29]  ( .D(data_out_b[29]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][29] ) );
  EDFFX1 \matrix_b_reg[4][29]  ( .D(data_out_b[29]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][29] ) );
  EDFFX1 \matrix_b_reg[3][29]  ( .D(data_out_b[29]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][29] ) );
  EDFFX1 \matrix_b_reg[0][28]  ( .D(data_out_b[28]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][28] ) );
  EDFFX1 \matrix_b_reg[8][28]  ( .D(data_out_b[28]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][28] ) );
  EDFFX1 \matrix_b_reg[6][28]  ( .D(data_out_b[28]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][28] ) );
  EDFFX1 \matrix_b_reg[5][28]  ( .D(data_out_b[28]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][28] ) );
  EDFFX1 \matrix_b_reg[4][28]  ( .D(data_out_b[28]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][28] ) );
  EDFFX1 \matrix_b_reg[3][28]  ( .D(data_out_b[28]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][28] ) );
  EDFFX1 \matrix_b_reg[0][27]  ( .D(data_out_b[27]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][27] ) );
  EDFFX1 \matrix_b_reg[8][27]  ( .D(data_out_b[27]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][27] ) );
  EDFFX1 \matrix_b_reg[6][27]  ( .D(data_out_b[27]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][27] ) );
  EDFFX1 \matrix_b_reg[5][27]  ( .D(data_out_b[27]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][27] ) );
  EDFFX1 \matrix_b_reg[4][27]  ( .D(data_out_b[27]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][27] ) );
  EDFFX1 \matrix_b_reg[3][27]  ( .D(data_out_b[27]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][27] ) );
  EDFFX1 \matrix_b_reg[0][26]  ( .D(data_out_b[26]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][26] ) );
  EDFFX1 \matrix_b_reg[8][26]  ( .D(data_out_b[26]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][26] ) );
  EDFFX1 \matrix_b_reg[6][26]  ( .D(data_out_b[26]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][26] ) );
  EDFFX1 \matrix_b_reg[5][26]  ( .D(data_out_b[26]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][26] ) );
  EDFFX1 \matrix_b_reg[4][26]  ( .D(data_out_b[26]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][26] ) );
  EDFFX1 \matrix_b_reg[3][26]  ( .D(data_out_b[26]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][26] ) );
  EDFFX1 \matrix_b_reg[0][25]  ( .D(data_out_b[25]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][25] ) );
  EDFFX1 \matrix_b_reg[8][25]  ( .D(data_out_b[25]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][25] ) );
  EDFFX1 \matrix_b_reg[6][25]  ( .D(data_out_b[25]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][25] ) );
  EDFFX1 \matrix_b_reg[5][25]  ( .D(data_out_b[25]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][25] ) );
  EDFFX1 \matrix_b_reg[4][25]  ( .D(data_out_b[25]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][25] ) );
  EDFFX1 \matrix_b_reg[3][25]  ( .D(data_out_b[25]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][25] ) );
  EDFFX1 \matrix_b_reg[0][24]  ( .D(data_out_b[24]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][24] ) );
  EDFFX1 \matrix_b_reg[8][24]  ( .D(data_out_b[24]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][24] ) );
  EDFFX1 \matrix_b_reg[6][24]  ( .D(data_out_b[24]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][24] ) );
  EDFFX1 \matrix_b_reg[5][24]  ( .D(data_out_b[24]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][24] ) );
  EDFFX1 \matrix_b_reg[4][24]  ( .D(data_out_b[24]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][24] ) );
  EDFFX1 \matrix_b_reg[3][24]  ( .D(data_out_b[24]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][24] ) );
  EDFFX1 \matrix_b_reg[7][23]  ( .D(data_out_b[23]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][23] ) );
  EDFFX1 \matrix_b_reg[0][23]  ( .D(data_out_b[23]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][23] ) );
  EDFFX1 \matrix_b_reg[8][23]  ( .D(data_out_b[23]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][23] ) );
  EDFFX1 \matrix_b_reg[6][23]  ( .D(data_out_b[23]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][23] ) );
  EDFFX1 \matrix_b_reg[2][23]  ( .D(data_out_b[23]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][23] ) );
  EDFFX1 \matrix_b_reg[3][23]  ( .D(data_out_b[23]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][23] ) );
  EDFFX1 \matrix_b_reg[7][22]  ( .D(data_out_b[22]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][22] ) );
  EDFFX1 \matrix_b_reg[0][22]  ( .D(data_out_b[22]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][22] ) );
  EDFFX1 \matrix_b_reg[8][22]  ( .D(data_out_b[22]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][22] ) );
  EDFFX1 \matrix_b_reg[6][22]  ( .D(data_out_b[22]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][22] ) );
  EDFFX1 \matrix_b_reg[2][22]  ( .D(data_out_b[22]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][22] ) );
  EDFFX1 \matrix_b_reg[3][22]  ( .D(data_out_b[22]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][22] ) );
  EDFFX1 \matrix_b_reg[7][21]  ( .D(data_out_b[21]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][21] ) );
  EDFFX1 \matrix_b_reg[0][21]  ( .D(data_out_b[21]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][21] ) );
  EDFFX1 \matrix_b_reg[8][21]  ( .D(data_out_b[21]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][21] ) );
  EDFFX1 \matrix_b_reg[6][21]  ( .D(data_out_b[21]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][21] ) );
  EDFFX1 \matrix_b_reg[2][21]  ( .D(data_out_b[21]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][21] ) );
  EDFFX1 \matrix_b_reg[3][21]  ( .D(data_out_b[21]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][21] ) );
  EDFFX1 \matrix_b_reg[8][20]  ( .D(data_out_b[20]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][20] ) );
  EDFFX1 \matrix_b_reg[7][20]  ( .D(data_out_b[20]), .E(n1570), .CK(clk), .Q(
        \matrix_b[7][20] ) );
  EDFFX1 \matrix_b_reg[0][20]  ( .D(data_out_b[20]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][20] ) );
  EDFFX1 \matrix_b_reg[6][20]  ( .D(data_out_b[20]), .E(n1556), .CK(clk), .Q(
        \matrix_b[6][20] ) );
  EDFFX1 \matrix_b_reg[2][20]  ( .D(data_out_b[20]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][20] ) );
  EDFFX1 \matrix_b_reg[3][20]  ( .D(data_out_b[20]), .E(n1908), .CK(clk), .Q(
        \matrix_b[3][20] ) );
  EDFFX1 \matrix_b_reg[8][15]  ( .D(data_out_b[15]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][15] ) );
  EDFFX1 \matrix_b_reg[0][15]  ( .D(data_out_b[15]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][15] ) );
  EDFFX1 \matrix_b_reg[5][15]  ( .D(data_out_b[15]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][15] ) );
  EDFFX1 \matrix_b_reg[2][15]  ( .D(data_out_b[15]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][15] ) );
  EDFFX1 \matrix_b_reg[1][15]  ( .D(data_out_b[15]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][15] ) );
  EDFFX1 \matrix_b_reg[8][14]  ( .D(data_out_b[14]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][14] ) );
  EDFFX1 \matrix_b_reg[0][14]  ( .D(data_out_b[14]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][14] ) );
  EDFFX1 \matrix_b_reg[5][14]  ( .D(data_out_b[14]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][14] ) );
  EDFFX1 \matrix_b_reg[2][14]  ( .D(data_out_b[14]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][14] ) );
  EDFFX1 \matrix_b_reg[1][14]  ( .D(data_out_b[14]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][14] ) );
  EDFFX1 \matrix_b_reg[8][13]  ( .D(data_out_b[13]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][13] ) );
  EDFFX1 \matrix_b_reg[0][13]  ( .D(data_out_b[13]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][13] ) );
  EDFFX1 \matrix_b_reg[5][13]  ( .D(data_out_b[13]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][13] ) );
  EDFFX1 \matrix_b_reg[2][13]  ( .D(data_out_b[13]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][13] ) );
  EDFFX1 \matrix_b_reg[1][13]  ( .D(data_out_b[13]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][13] ) );
  EDFFX1 \matrix_b_reg[0][12]  ( .D(data_out_b[12]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][12] ) );
  EDFFX1 \matrix_b_reg[8][12]  ( .D(data_out_b[12]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][12] ) );
  EDFFX1 \matrix_b_reg[5][12]  ( .D(data_out_b[12]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][12] ) );
  EDFFX1 \matrix_b_reg[2][12]  ( .D(data_out_b[12]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][12] ) );
  EDFFX1 \matrix_b_reg[1][12]  ( .D(data_out_b[12]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][12] ) );
  EDFFX1 \matrix_b_reg[0][11]  ( .D(data_out_b[11]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][11] ) );
  EDFFX1 \matrix_b_reg[8][11]  ( .D(data_out_b[11]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][11] ) );
  EDFFX1 \matrix_b_reg[5][11]  ( .D(data_out_b[11]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][11] ) );
  EDFFX1 \matrix_b_reg[2][11]  ( .D(data_out_b[11]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][11] ) );
  EDFFX1 \matrix_b_reg[1][11]  ( .D(data_out_b[11]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][11] ) );
  EDFFX1 \matrix_b_reg[0][10]  ( .D(data_out_b[10]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][10] ) );
  EDFFX1 \matrix_b_reg[8][10]  ( .D(data_out_b[10]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][10] ) );
  EDFFX1 \matrix_b_reg[5][10]  ( .D(data_out_b[10]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][10] ) );
  EDFFX1 \matrix_b_reg[2][10]  ( .D(data_out_b[10]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][10] ) );
  EDFFX1 \matrix_b_reg[1][10]  ( .D(data_out_b[10]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][10] ) );
  EDFFX1 \matrix_b_reg[0][9]  ( .D(data_out_b[9]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][9] ) );
  EDFFX1 \matrix_b_reg[8][9]  ( .D(data_out_b[9]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][9] ) );
  EDFFX1 \matrix_b_reg[5][9]  ( .D(data_out_b[9]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][9] ) );
  EDFFX1 \matrix_b_reg[2][9]  ( .D(data_out_b[9]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][9] ) );
  EDFFX1 \matrix_b_reg[1][9]  ( .D(data_out_b[9]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][9] ) );
  EDFFX1 \matrix_b_reg[0][8]  ( .D(data_out_b[8]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][8] ) );
  EDFFX1 \matrix_b_reg[8][8]  ( .D(data_out_b[8]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][8] ) );
  EDFFX1 \matrix_b_reg[5][8]  ( .D(data_out_b[8]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][8] ) );
  EDFFX1 \matrix_b_reg[2][8]  ( .D(data_out_b[8]), .E(n1558), .CK(clk), .Q(
        \matrix_b[2][8] ) );
  EDFFX1 \matrix_b_reg[1][8]  ( .D(data_out_b[8]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][8] ) );
  EDFFX1 \matrix_b_reg[0][7]  ( .D(data_out_b[7]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][7] ) );
  EDFFX1 \matrix_b_reg[8][7]  ( .D(data_out_b[7]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][7] ) );
  EDFFX1 \matrix_b_reg[5][7]  ( .D(data_out_b[7]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][7] ) );
  EDFFX1 \matrix_b_reg[4][7]  ( .D(data_out_b[7]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][7] ) );
  EDFFX1 \matrix_b_reg[1][7]  ( .D(data_out_b[7]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][7] ) );
  EDFFX1 \matrix_b_reg[0][6]  ( .D(data_out_b[6]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][6] ) );
  EDFFX1 \matrix_b_reg[8][6]  ( .D(data_out_b[6]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][6] ) );
  EDFFX1 \matrix_b_reg[5][6]  ( .D(data_out_b[6]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][6] ) );
  EDFFX1 \matrix_b_reg[4][6]  ( .D(data_out_b[6]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][6] ) );
  EDFFX1 \matrix_b_reg[1][6]  ( .D(data_out_b[6]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][6] ) );
  EDFFX1 \matrix_b_reg[0][5]  ( .D(data_out_b[5]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][5] ) );
  EDFFX1 \matrix_b_reg[8][5]  ( .D(data_out_b[5]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][5] ) );
  EDFFX1 \matrix_b_reg[5][5]  ( .D(data_out_b[5]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][5] ) );
  EDFFX1 \matrix_b_reg[4][5]  ( .D(data_out_b[5]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][5] ) );
  EDFFX1 \matrix_b_reg[1][5]  ( .D(data_out_b[5]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][5] ) );
  EDFFX1 \matrix_b_reg[0][4]  ( .D(data_out_b[4]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][4] ) );
  EDFFX1 \matrix_b_reg[8][4]  ( .D(data_out_b[4]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][4] ) );
  EDFFX1 \matrix_b_reg[5][4]  ( .D(data_out_b[4]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][4] ) );
  EDFFX1 \matrix_b_reg[4][4]  ( .D(data_out_b[4]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][4] ) );
  EDFFX1 \matrix_b_reg[1][4]  ( .D(data_out_b[4]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][4] ) );
  EDFFX1 \matrix_b_reg[0][3]  ( .D(data_out_b[3]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][3] ) );
  EDFFX1 \matrix_b_reg[8][3]  ( .D(data_out_b[3]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][3] ) );
  EDFFX1 \matrix_b_reg[5][3]  ( .D(data_out_b[3]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][3] ) );
  EDFFX1 \matrix_b_reg[4][3]  ( .D(data_out_b[3]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][3] ) );
  EDFFX1 \matrix_b_reg[1][3]  ( .D(data_out_b[3]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][3] ) );
  EDFFX1 \matrix_b_reg[0][2]  ( .D(data_out_b[2]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][2] ) );
  EDFFX1 \matrix_b_reg[8][2]  ( .D(data_out_b[2]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][2] ) );
  EDFFX1 \matrix_b_reg[5][2]  ( .D(data_out_b[2]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][2] ) );
  EDFFX1 \matrix_b_reg[4][2]  ( .D(data_out_b[2]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][2] ) );
  EDFFX1 \matrix_b_reg[1][2]  ( .D(data_out_b[2]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][2] ) );
  EDFFX1 \matrix_b_reg[0][1]  ( .D(data_out_b[1]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][1] ) );
  EDFFX1 \matrix_b_reg[8][1]  ( .D(data_out_b[1]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][1] ) );
  EDFFX1 \matrix_b_reg[5][1]  ( .D(data_out_b[1]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][1] ) );
  EDFFX1 \matrix_b_reg[4][1]  ( .D(data_out_b[1]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][1] ) );
  EDFFX1 \matrix_b_reg[1][1]  ( .D(data_out_b[1]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][1] ) );
  EDFFX1 \matrix_b_reg[0][0]  ( .D(data_out_b[0]), .E(n1546), .CK(clk), .Q(
        \matrix_b[0][0] ) );
  EDFFX1 \matrix_b_reg[8][0]  ( .D(data_out_b[0]), .E(n1561), .CK(clk), .Q(
        \matrix_b[8][0] ) );
  EDFFX1 \matrix_b_reg[5][0]  ( .D(data_out_b[0]), .E(n1563), .CK(clk), .Q(
        \matrix_b[5][0] ) );
  EDFFX1 \matrix_b_reg[4][0]  ( .D(data_out_b[0]), .E(n1564), .CK(clk), .Q(
        \matrix_b[4][0] ) );
  EDFFX1 \matrix_b_reg[1][0]  ( .D(data_out_b[0]), .E(n1567), .CK(clk), .Q(
        \matrix_b[1][0] ) );
  DFFQX1 wr_en_out_reg ( .D(n1499), .CK(clk), .Q(wr_en_out) );
  ADDHXL \add_332/U1_1_3  ( .A(k[3]), .B(\add_332/carry[3] ), .CO(N722), .S(
        N721) );
  ADDFHX2 \add_357/U1_3  ( .A(k[3]), .B(n[3]), .CI(\add_357/carry[3] ), .CO(
        N783), .S(N782) );
  ADDFX2 \add_357_2/U1_2  ( .A(N247), .B(n[1]), .CI(n1518), .CO(
        \add_357_2/carry[3] ), .S(N787) );
  AOI221X1 U1000 ( .A0(n1628), .A1(n1717), .B0(n1712), .B1(n1711), .C0(n1710), 
        .Y(n1713) );
  BUFX4 U1001 ( .A(n876), .Y(n1615) );
  NAND2XL U1002 ( .A(n1753), .B(n1614), .Y(n876) );
  AND2X4 U1003 ( .A(n820), .B(n808), .Y(n822) );
  NOR2X4 U1004 ( .A(n1540), .B(n807), .Y(n808) );
  BUFX4 U1005 ( .A(n877), .Y(n1616) );
  OAI222X4 U1006 ( .A0(n1615), .A1(n704), .B0(n1758), .B1(n877), .C0(n1542), 
        .C1(n736), .Y(n1326) );
  OAI222X4 U1007 ( .A0(n1615), .A1(n706), .B0(n1760), .B1(n877), .C0(n1542), 
        .C1(n738), .Y(n1328) );
  OAI222X4 U1008 ( .A0(n1615), .A1(n708), .B0(n1762), .B1(n877), .C0(n1542), 
        .C1(n740), .Y(n1330) );
  OAI222X4 U1009 ( .A0(n1615), .A1(n703), .B0(n1757), .B1(n877), .C0(n1542), 
        .C1(n735), .Y(n1325) );
  OAI222X4 U1010 ( .A0(n1615), .A1(n705), .B0(n1759), .B1(n877), .C0(n1542), 
        .C1(n737), .Y(n1327) );
  NAND2X2 U1011 ( .A(n906), .B(n1614), .Y(n877) );
  NOR2X6 U1012 ( .A(n1528), .B(n1529), .Y(n1543) );
  INVX3 U1013 ( .A(n[0]), .Y(n1528) );
  CLKINVX1 U1014 ( .A(N787), .Y(n1744) );
  INVX4 U1015 ( .A(n1618), .Y(n1752) );
  BUFX4 U1016 ( .A(n905), .Y(n1617) );
  INVX4 U1017 ( .A(n1544), .Y(n1540) );
  AO21X1 U1018 ( .A0(n1743), .A1(n1732), .B0(N786), .Y(n1731) );
  CLKINVX1 U1019 ( .A(n911), .Y(n1753) );
  OAI211X1 U1020 ( .A0(n912), .A1(n913), .B0(n910), .C0(n909), .Y(n911) );
  NAND3X1 U1021 ( .A(n914), .B(n915), .C(n916), .Y(n913) );
  INVX8 U1022 ( .A(N785), .Y(n1529) );
  OAI21XL U1023 ( .A0(n819), .A1(n1855), .B0(n1854), .Y(n1278) );
  CLKINVX1 U1024 ( .A(rst), .Y(n1520) );
  OA21XL U1025 ( .A0(n1282), .A1(n1854), .B0(n1278), .Y(n1276) );
  NOR2BX2 U1026 ( .AN(n1545), .B(n941), .Y(n907) );
  OR4X1 U1027 ( .A(n1626), .B(n1621), .C(n1727), .D(n1726), .Y(n1545) );
  NAND2X1 U1028 ( .A(n1526), .B(n784), .Y(n1499) );
  AND2X2 U1029 ( .A(data_in_o[18]), .B(n1540), .Y(n1541) );
  NAND2X1 U1030 ( .A(n822), .B(n827), .Y(n1523) );
  NAND2X1 U1031 ( .A(temp1[18]), .B(n1752), .Y(n1524) );
  AND2X2 U1032 ( .A(data_in_o[20]), .B(n797), .Y(n1534) );
  AND2X2 U1033 ( .A(data_in_o[21]), .B(n797), .Y(n1530) );
  OAI22XL U1034 ( .A0(n1714), .A1(n1713), .B0(N783), .B1(n1533), .Y(n1716) );
  OAI21X1 U1035 ( .A0(n819), .A1(n807), .B0(n1544), .Y(n838) );
  AND3X2 U1036 ( .A(n1690), .B(n1692), .C(n1146), .Y(n1510) );
  INVXL U1037 ( .A(index_a[2]), .Y(n1693) );
  CLKINVX3 U1038 ( .A(n1544), .Y(n797) );
  OR3X2 U1039 ( .A(n1548), .B(n1549), .C(n1550), .Y(n1511) );
  OR3X2 U1040 ( .A(n1537), .B(n1538), .C(n1539), .Y(n1512) );
  OR3X2 U1041 ( .A(n1534), .B(n1535), .C(n1536), .Y(n1513) );
  OR3X2 U1042 ( .A(n1530), .B(n1531), .C(n1532), .Y(n1514) );
  AND3X2 U1043 ( .A(n909), .B(n910), .C(n907), .Y(n1562) );
  AND2X2 U1044 ( .A(N785), .B(n[0]), .Y(n1517) );
  AND3X4 U1045 ( .A(N784), .B(n1906), .C(N791), .Y(n1544) );
  AND2X2 U1046 ( .A(n[0]), .B(N241), .Y(n1518) );
  CLKINVX1 U1047 ( .A(n971), .Y(n1653) );
  CLKINVX1 U1048 ( .A(n972), .Y(n1650) );
  INVX6 U1049 ( .A(n1520), .Y(n1521) );
  CLKAND2X3 U1050 ( .A(n1058), .B(n1690), .Y(n1568) );
  AND3X4 U1051 ( .A(n1683), .B(n1681), .C(n1268), .Y(n1556) );
  INVX3 U1052 ( .A(n1594), .Y(n1908) );
  AND3X6 U1053 ( .A(n1691), .B(n1690), .C(n1146), .Y(n1565) );
  AND3X6 U1054 ( .A(n1689), .B(n1692), .C(n1146), .Y(n1566) );
  CLKAND2X6 U1055 ( .A(n1058), .B(n1689), .Y(n1559) );
  CLKAND2X6 U1056 ( .A(n1681), .B(n1274), .Y(n1561) );
  AND4XL U1057 ( .A(n1687), .B(n1272), .C(n1275), .D(n1907), .Y(n1274) );
  AND3X6 U1058 ( .A(n1683), .B(n1682), .C(n1268), .Y(n1563) );
  AND3X6 U1059 ( .A(n1681), .B(n1684), .C(n1268), .Y(n1564) );
  CLKAND2X6 U1060 ( .A(n1224), .B(n1682), .Y(n1567) );
  NOR3BX1 U1061 ( .AN(n1198), .B(n1684), .C(n1685), .Y(n1224) );
  CLKAND2X6 U1062 ( .A(n1151), .B(n1690), .Y(n1569) );
  AND4XL U1063 ( .A(n788), .B(n1694), .C(n1153), .D(n1907), .Y(n1151) );
  CLKAND2X6 U1064 ( .A(n1224), .B(n1681), .Y(n1558) );
  AND4X6 U1065 ( .A(n1198), .B(n1681), .C(n1684), .D(n1686), .Y(n1546) );
  AND4X6 U1066 ( .A(n1014), .B(n1689), .C(n1692), .D(n1693), .Y(n1547) );
  CLKAND2X6 U1067 ( .A(n1151), .B(n1689), .Y(n1560) );
  CLKAND2X6 U1068 ( .A(n1274), .B(n1682), .Y(n1570) );
  NOR4X4 U1069 ( .A(n1703), .B(n1702), .C(n1627), .D(n1628), .Y(N894) );
  NOR4BBX4 U1070 ( .AN(n1706), .BN(n1705), .C(n1625), .D(n1626), .Y(N892) );
  NOR4BBX4 U1071 ( .AN(n1700), .BN(n1699), .C(n1625), .D(n1626), .Y(N896) );
  NAND3BX1 U1072 ( .AN(n1541), .B(n1523), .C(n1524), .Y(n1522) );
  OAI22X1 U1073 ( .A0(n1708), .A1(n1515), .B0(N782), .B1(n1708), .Y(n1711) );
  NAND2X1 U1074 ( .A(N247), .B(\add_357/carry[2] ), .Y(n1553) );
  AOI221X1 U1075 ( .A0(n1628), .A1(n1728), .B0(n1723), .B1(n1722), .C0(n1721), 
        .Y(n1724) );
  OAI22X1 U1076 ( .A0(n1719), .A1(n1515), .B0(N714), .B1(n1719), .Y(n1722) );
  NOR2X1 U1077 ( .A(n807), .B(n805), .Y(n1525) );
  OR2X4 U1078 ( .A(n1525), .B(n797), .Y(n810) );
  INVX3 U1079 ( .A(n1540), .Y(n1680) );
  OAI221X1 U1080 ( .A0(n1772), .A1(n809), .B0(n810), .B1(n710), .C0(n817), .Y(
        n1297) );
  OAI221X1 U1081 ( .A0(n1774), .A1(n809), .B0(n810), .B1(n712), .C0(n815), .Y(
        n1295) );
  OAI221X1 U1082 ( .A0(n1776), .A1(n809), .B0(n810), .B1(n714), .C0(n813), .Y(
        n1293) );
  OAI221X1 U1083 ( .A0(n1778), .A1(n809), .B0(n810), .B1(n716), .C0(n811), .Y(
        n1291) );
  OAI221X1 U1084 ( .A0(n1771), .A1(n809), .B0(n810), .B1(n709), .C0(n818), .Y(
        n1298) );
  OAI221X1 U1085 ( .A0(n1773), .A1(n809), .B0(n810), .B1(n711), .C0(n816), .Y(
        n1296) );
  OAI221X1 U1086 ( .A0(n1775), .A1(n809), .B0(n810), .B1(n713), .C0(n814), .Y(
        n1294) );
  OAI221X1 U1087 ( .A0(n1777), .A1(n809), .B0(n810), .B1(n715), .C0(n812), .Y(
        n1292) );
  OR3X2 U1088 ( .A(n1748), .B(n783), .C(n1754), .Y(n1526) );
  AND2X2 U1089 ( .A(n1906), .B(N793), .Y(n1527) );
  NOR2X1 U1090 ( .A(n1527), .B(n1680), .Y(n783) );
  INVXL U1091 ( .A(N791), .Y(n1748) );
  INVXL U1092 ( .A(N784), .Y(n1754) );
  AND2XL U1093 ( .A(n822), .B(n833), .Y(n1531) );
  AND2XL U1094 ( .A(temp1[21]), .B(n1752), .Y(n1532) );
  OR4X2 U1095 ( .A(n1626), .B(n1621), .C(n1716), .D(n1715), .Y(N784) );
  AND2XL U1096 ( .A(n822), .B(n831), .Y(n1535) );
  AND2XL U1097 ( .A(temp1[20]), .B(n1752), .Y(n1536) );
  CLKINVX1 U1098 ( .A(n1573), .Y(n1747) );
  AND2XL U1099 ( .A(temp1[16]), .B(n1752), .Y(n1539) );
  AND2X1 U1100 ( .A(n822), .B(n823), .Y(n1538) );
  AOI222X1 U1101 ( .A0(data_in_o[19]), .A1(n797), .B0(n822), .B1(n829), .C0(
        temp1[19]), .C1(n1752), .Y(n828) );
  AOI222X1 U1102 ( .A0(data_in_o[22]), .A1(n797), .B0(n822), .B1(n835), .C0(
        temp1[22]), .C1(n1752), .Y(n834) );
  AOI222X1 U1103 ( .A0(data_in_o[23]), .A1(n797), .B0(n822), .B1(n837), .C0(
        temp1[23]), .C1(n1752), .Y(n836) );
  INVX3 U1104 ( .A(N789), .Y(n1746) );
  AND2XL U1105 ( .A(data_in_o[16]), .B(n797), .Y(n1537) );
  OAI211X1 U1106 ( .A0(n1792), .A1(n1674), .B0(n870), .C0(n871), .Y(n827) );
  XOR2X1 U1107 ( .A(k[3]), .B(n1574), .Y(N733) );
  XOR2X1 U1108 ( .A(k[3]), .B(n1575), .Y(N727) );
  XOR2X1 U1109 ( .A(\add_357/carry[2] ), .B(n1551), .Y(N781) );
  CLKBUFX3 U1110 ( .A(n1614), .Y(n1542) );
  BUFX6 U1111 ( .A(n878), .Y(n1614) );
  OAI22XL U1112 ( .A0(N782), .A1(n1515), .B0(N782), .B1(n1709), .Y(n1710) );
  OAI22X1 U1113 ( .A0(N714), .A1(n1515), .B0(N714), .B1(n1720), .Y(n1721) );
  INVX1 U1114 ( .A(n1720), .Y(n1728) );
  NAND3X2 U1115 ( .A(n1552), .B(n1553), .C(n1554), .Y(\add_357/carry[3] ) );
  NAND2X1 U1116 ( .A(n1628), .B(n1745), .Y(n1735) );
  NOR2X2 U1117 ( .A(n909), .B(n1852), .Y(n906) );
  AND2X2 U1118 ( .A(n1697), .B(n1696), .Y(N898) );
  AND2XL U1119 ( .A(temp1[17]), .B(n1752), .Y(n1550) );
  NAND3X2 U1120 ( .A(N785), .B(n1856), .C(n808), .Y(n794) );
  NAND4X4 U1121 ( .A(n942), .B(n918), .C(n943), .D(n944), .Y(n910) );
  OAI31X4 U1122 ( .A0(n805), .A1(n806), .A2(n807), .B0(n1680), .Y(n795) );
  INVXL U1123 ( .A(n1709), .Y(n1717) );
  OAI221X1 U1124 ( .A0(n1629), .A1(n1744), .B0(n1628), .B1(n1745), .C0(n1733), 
        .Y(n1734) );
  OAI211XL U1125 ( .A0(n1732), .A1(n1743), .B0(n1731), .C0(n1730), .Y(n1733)
         );
  NAND4XL U1126 ( .A(n1735), .B(n1730), .C(n1516), .D(n1519), .Y(n1742) );
  NAND2X1 U1127 ( .A(n1855), .B(n1854), .Y(n807) );
  CLKBUFX3 U1128 ( .A(n970), .Y(n1595) );
  CLKBUFX3 U1129 ( .A(n975), .Y(n1604) );
  CLKINVX1 U1130 ( .A(n972), .Y(n1651) );
  INVX3 U1131 ( .A(n1690), .Y(n1689) );
  CLKINVX1 U1132 ( .A(n1684), .Y(n1683) );
  INVX3 U1133 ( .A(n1682), .Y(n1681) );
  NOR3BXL U1134 ( .AN(n1014), .B(n1692), .C(index_a[2]), .Y(n1058) );
  CLKINVX1 U1135 ( .A(n1686), .Y(n1685) );
  NAND2XL U1136 ( .A(wr_en_out), .B(n783), .Y(n784) );
  NOR3X2 U1137 ( .A(n945), .B(n946), .C(n947), .Y(n944) );
  XOR2XL U1138 ( .A(n[0]), .B(N241), .Y(N786) );
  XNOR2XL U1139 ( .A(N241), .B(N785), .Y(N731) );
  XOR2XL U1140 ( .A(N247), .B(\add_332_3/carry[2] ), .Y(N732) );
  XNOR2XL U1141 ( .A(n1630), .B(N241), .Y(n953) );
  XOR2XL U1142 ( .A(counter[0]), .B(N785), .Y(n915) );
  XOR2XL U1143 ( .A(N247), .B(N241), .Y(N726) );
  OR2XL U1144 ( .A(N241), .B(N785), .Y(\add_332_3/carry[2] ) );
  XOR2XL U1145 ( .A(N785), .B(n[0]), .Y(N794) );
  NAND2XL U1146 ( .A(k[3]), .B(n1574), .Y(n1577) );
  AND2XL U1147 ( .A(N247), .B(\add_332_3/carry[2] ), .Y(n1574) );
  AND2XL U1148 ( .A(N247), .B(N241), .Y(n1575) );
  AND2XL U1149 ( .A(k[3]), .B(n1575), .Y(n1576) );
  CLKBUFX3 U1150 ( .A(counter[2]), .Y(n1629) );
  BUFX4 U1151 ( .A(counter[3]), .Y(n1628) );
  INVX1 U1152 ( .A(k[3]), .Y(n1854) );
  INVX1 U1153 ( .A(N247), .Y(n1855) );
  NOR2XL U1154 ( .A(n1856), .B(N785), .Y(n806) );
  AOI22XL U1155 ( .A0(N247), .A1(n1277), .B0(n1855), .B1(n1276), .Y(n1279) );
  NOR2BXL U1156 ( .AN(n819), .B(N247), .Y(n1282) );
  INVX1 U1157 ( .A(N241), .Y(n1856) );
  NOR2X1 U1158 ( .A(N785), .B(N241), .Y(n819) );
  XOR2XL U1159 ( .A(k[3]), .B(n1694), .Y(n791) );
  XOR2XL U1160 ( .A(N241), .B(n1691), .Y(n792) );
  NAND2BXL U1161 ( .AN(k[3]), .B(n1855), .Y(\sub_142/carry[4] ) );
  XNOR2XL U1162 ( .A(k[3]), .B(N247), .Y(N243) );
  NOR2X1 U1163 ( .A(n700), .B(n1629), .Y(n1197) );
  NOR2X1 U1164 ( .A(n699), .B(n1628), .Y(n1225) );
  NAND2X1 U1165 ( .A(cur_state[0]), .B(n163), .Y(n785) );
  NOR4X1 U1166 ( .A(n1695), .B(index_a[5]), .C(index_a[6]), .D(index_a[7]), 
        .Y(n788) );
  CLKINVX1 U1167 ( .A(index_a[0]), .Y(n1690) );
  CLKINVX1 U1168 ( .A(index_a[1]), .Y(n1692) );
  CLKINVX1 U1169 ( .A(index_b[0]), .Y(n1682) );
  CLKINVX1 U1170 ( .A(index_b[1]), .Y(n1684) );
  CLKINVX1 U1171 ( .A(index_b[2]), .Y(n1686) );
  AND4X1 U1172 ( .A(l[1]), .B(l[0]), .C(n957), .D(n629), .Y(n844) );
  AND4X1 U1173 ( .A(l[0]), .B(n957), .C(n630), .D(n629), .Y(n841) );
  AND4X1 U1174 ( .A(l[1]), .B(n957), .C(n631), .D(n629), .Y(n840) );
  XOR2X1 U1175 ( .A(n[2]), .B(N247), .Y(n1551) );
  NAND2XL U1176 ( .A(n[2]), .B(\add_357/carry[2] ), .Y(n1552) );
  NAND2XL U1177 ( .A(N247), .B(n[2]), .Y(n1554) );
  AND2X2 U1178 ( .A(data_in_o[17]), .B(n1540), .Y(n1548) );
  AND2XL U1179 ( .A(n822), .B(n825), .Y(n1549) );
  CLKBUFX3 U1180 ( .A(n1205), .Y(n1640) );
  CLKBUFX3 U1181 ( .A(n1206), .Y(n1639) );
  NOR2X1 U1182 ( .A(n1641), .B(n1664), .Y(n1206) );
  NOR2X1 U1183 ( .A(n1641), .B(n1662), .Y(n1205) );
  INVX3 U1184 ( .A(n1510), .Y(n1645) );
  INVX3 U1185 ( .A(n1510), .Y(n1646) );
  CLKBUFX3 U1186 ( .A(n1215), .Y(n1638) );
  CLKBUFX3 U1187 ( .A(n1216), .Y(n1637) );
  NAND2X2 U1188 ( .A(n1605), .B(n1668), .Y(n1199) );
  NAND2X2 U1189 ( .A(n1605), .B(n1909), .Y(n1200) );
  NAND2X2 U1190 ( .A(n1597), .B(n1911), .Y(n1264) );
  INVX3 U1191 ( .A(n973), .Y(n1912) );
  NOR2X1 U1192 ( .A(n1643), .B(n1670), .Y(n1216) );
  NOR2X1 U1193 ( .A(n1643), .B(n1659), .Y(n1215) );
  NAND4X1 U1194 ( .A(n1139), .B(n1140), .C(n1656), .D(n965), .Y(n1052) );
  NOR2X1 U1195 ( .A(n1571), .B(n1663), .Y(n1140) );
  CLKBUFX3 U1196 ( .A(n1163), .Y(n1643) );
  CLKBUFX3 U1197 ( .A(n1196), .Y(n1641) );
  CLKBUFX3 U1198 ( .A(n1016), .Y(n1612) );
  NAND2X1 U1199 ( .A(n1857), .B(n1008), .Y(n1016) );
  CLKBUFX3 U1200 ( .A(n1908), .Y(n1634) );
  INVX3 U1201 ( .A(n1571), .Y(n1664) );
  INVX3 U1202 ( .A(n1663), .Y(n1662) );
  INVX3 U1203 ( .A(n1571), .Y(n1665) );
  INVX3 U1204 ( .A(n1668), .Y(n1666) );
  CLKBUFX3 U1205 ( .A(n1243), .Y(n1599) );
  NAND2X1 U1206 ( .A(n1598), .B(n1668), .Y(n1243) );
  CLKBUFX3 U1207 ( .A(n1203), .Y(n1603) );
  NAND2X1 U1208 ( .A(n1601), .B(n1653), .Y(n1203) );
  CLKBUFX3 U1209 ( .A(n1510), .Y(n1647) );
  CLKBUFX3 U1210 ( .A(n1510), .Y(n1648) );
  INVX3 U1211 ( .A(n1653), .Y(n1652) );
  CLKBUFX3 U1212 ( .A(n1163), .Y(n1644) );
  CLKBUFX3 U1213 ( .A(n1196), .Y(n1642) );
  CLKBUFX3 U1214 ( .A(n1556), .Y(n1633) );
  CLKBUFX3 U1215 ( .A(n1557), .Y(n1635) );
  CLKINVX1 U1216 ( .A(n1668), .Y(n1667) );
  OA21XL U1217 ( .A0(n1754), .A1(n1748), .B0(N793), .Y(n1555) );
  OAI21X2 U1218 ( .A0(n906), .A1(n1852), .B0(n1617), .Y(n904) );
  NAND2X2 U1219 ( .A(n1617), .B(n1753), .Y(n903) );
  OA21XL U1220 ( .A0(n906), .A1(n1753), .B0(n907), .Y(n878) );
  NOR2BX1 U1221 ( .AN(n907), .B(n908), .Y(n905) );
  AOI211X1 U1222 ( .A0(n1853), .A1(n906), .B0(n1753), .C0(n1852), .Y(n908) );
  CLKINVX1 U1223 ( .A(n807), .Y(n1853) );
  CLKBUFX3 U1224 ( .A(n1562), .Y(n1632) );
  AO22X1 U1225 ( .A0(n1689), .A1(n1619), .B0(N257), .B1(n1620), .Y(n1506) );
  AO22X1 U1226 ( .A0(n1681), .A1(n1619), .B0(N265), .B1(n1620), .Y(n1497) );
  AO22X1 U1227 ( .A0(index_a[2]), .A1(n1619), .B0(N259), .B1(n1620), .Y(n1504)
         );
  AO22X1 U1228 ( .A0(n1691), .A1(n1619), .B0(N258), .B1(n1620), .Y(n1505) );
  AO22X1 U1229 ( .A0(n1619), .A1(n1685), .B0(N267), .B1(n1620), .Y(n1495) );
  AO22X1 U1230 ( .A0(n1619), .A1(n1683), .B0(N266), .B1(n1620), .Y(n1496) );
  NAND2X2 U1231 ( .A(n1597), .B(n1657), .Y(n1263) );
  NAND2X2 U1232 ( .A(n1164), .B(n1165), .Y(n973) );
  NAND3BX1 U1233 ( .AN(n1052), .B(n1604), .C(n1652), .Y(n1008) );
  AND3X2 U1234 ( .A(n1691), .B(n1689), .C(n1146), .Y(n1557) );
  CLKBUFX3 U1235 ( .A(n1186), .Y(n1601) );
  AOI2BB1X1 U1236 ( .A0N(n1654), .A1N(n1657), .B0(n1596), .Y(n1186) );
  NOR2X1 U1237 ( .A(n1671), .B(n1660), .Y(n1139) );
  CLKINVX1 U1238 ( .A(n1596), .Y(n1857) );
  INVX3 U1239 ( .A(n974), .Y(n1910) );
  CLKBUFX3 U1240 ( .A(n1245), .Y(n1598) );
  AOI2BB1X1 U1241 ( .A0N(n1651), .A1N(n1668), .B0(n1596), .Y(n1245) );
  CLKBUFX3 U1242 ( .A(n1177), .Y(n1607) );
  AOI2BB1X1 U1243 ( .A0N(n1596), .A1N(n1595), .B0(n1601), .Y(n1177) );
  CLKBUFX3 U1244 ( .A(n1167), .Y(n1608) );
  AOI2BB1X1 U1245 ( .A0N(n1596), .A1N(n1649), .B0(n1605), .Y(n1167) );
  CLKBUFX3 U1246 ( .A(n1154), .Y(n1609) );
  OA21XL U1247 ( .A0(n1596), .A1(n973), .B0(n1644), .Y(n1154) );
  CLKBUFX3 U1248 ( .A(n1187), .Y(n1606) );
  OA21XL U1249 ( .A0(n1596), .A1(n974), .B0(n1642), .Y(n1187) );
  CLKBUFX3 U1250 ( .A(n959), .Y(n1613) );
  OAI31XL U1251 ( .A0(n1007), .A1(n1910), .A2(n1008), .B0(n1857), .Y(n959) );
  NAND3X1 U1252 ( .A(n1649), .B(n973), .C(n1595), .Y(n1007) );
  CLKBUFX3 U1253 ( .A(n1060), .Y(n1611) );
  OAI31XL U1254 ( .A0(n1052), .A1(n1650), .A2(n1653), .B0(n1857), .Y(n1060) );
  CLKBUFX3 U1255 ( .A(n1102), .Y(n1610) );
  OAI31XL U1256 ( .A0(n1052), .A1(n1650), .A2(n1911), .B0(n1857), .Y(n1102) );
  INVX3 U1257 ( .A(n1650), .Y(n1649) );
  INVX3 U1258 ( .A(n1671), .Y(n1670) );
  INVX3 U1259 ( .A(n1660), .Y(n1658) );
  OR2X1 U1260 ( .A(n1139), .B(n1596), .Y(n1163) );
  OR2X1 U1261 ( .A(n1140), .B(n1596), .Y(n1196) );
  CLKBUFX3 U1262 ( .A(n1202), .Y(n1602) );
  NAND2X1 U1263 ( .A(n1601), .B(n1657), .Y(n1202) );
  CLKBUFX3 U1264 ( .A(n1244), .Y(n1600) );
  NAND2X1 U1265 ( .A(n1598), .B(n1650), .Y(n1244) );
  INVX3 U1266 ( .A(n1657), .Y(n1656) );
  CLKBUFX3 U1267 ( .A(n1176), .Y(n1605) );
  AOI2BB1X1 U1268 ( .A0N(n1909), .A1N(n1668), .B0(n1596), .Y(n1176) );
  INVX3 U1269 ( .A(n1595), .Y(n1911) );
  CLKBUFX3 U1270 ( .A(n1265), .Y(n1597) );
  AOI2BB1X1 U1271 ( .A0N(n1911), .A1N(n1657), .B0(n1596), .Y(n1265) );
  CLKBUFX3 U1272 ( .A(n1568), .Y(n1636) );
  INVX3 U1273 ( .A(n1604), .Y(n1909) );
  INVX3 U1274 ( .A(n965), .Y(n1668) );
  CLKINVX1 U1275 ( .A(n971), .Y(n1654) );
  CLKINVX1 U1276 ( .A(n1660), .Y(n1659) );
  INVX3 U1277 ( .A(n1661), .Y(n1663) );
  NAND2X2 U1278 ( .A(n806), .B(n808), .Y(n809) );
  CLKBUFX3 U1279 ( .A(n838), .Y(n1618) );
  CLKINVX1 U1280 ( .A(N788), .Y(n1745) );
  XOR2X1 U1281 ( .A(n1628), .B(N721), .Y(n945) );
  XOR2X1 U1282 ( .A(n1630), .B(N719), .Y(n947) );
  XOR2X1 U1283 ( .A(n1629), .B(N720), .Y(n946) );
  NAND3X1 U1284 ( .A(n917), .B(n918), .C(n919), .Y(n912) );
  CLKINVX1 U1285 ( .A(n910), .Y(n1852) );
  NOR2XL U1286 ( .A(N896), .B(n1794), .Y(psum3[0]) );
  NOR2XL U1287 ( .A(N892), .B(n1770), .Y(psum1[0]) );
  NOR2XL U1288 ( .A(N894), .B(n1786), .Y(psum2[0]) );
  NOR2X1 U1289 ( .A(n1854), .B(n1282), .Y(n1277) );
  NAND4X1 U1290 ( .A(n787), .B(n788), .C(n789), .D(n790), .Y(n786) );
  NOR2X1 U1291 ( .A(n791), .B(n792), .Y(n790) );
  XOR2X1 U1292 ( .A(n1529), .B(n1689), .Y(n787) );
  XOR2X1 U1293 ( .A(n1855), .B(index_a[2]), .Y(n789) );
  NOR2X1 U1294 ( .A(n1856), .B(n1529), .Y(n820) );
  CLKBUFX3 U1295 ( .A(n782), .Y(n1620) );
  NOR2BX1 U1296 ( .AN(n786), .B(n785), .Y(n782) );
  OR2X1 U1297 ( .A(n819), .B(n820), .Y(n805) );
  NOR2XL U1298 ( .A(N894), .B(n1784), .Y(psum2[2]) );
  NOR2XL U1299 ( .A(N894), .B(n1783), .Y(psum2[3]) );
  NOR2XL U1300 ( .A(N894), .B(n1782), .Y(psum2[4]) );
  NOR2XL U1301 ( .A(N894), .B(n1781), .Y(psum2[5]) );
  NOR2XL U1302 ( .A(N894), .B(n1780), .Y(psum2[6]) );
  NOR2XL U1303 ( .A(N896), .B(n1793), .Y(psum3[1]) );
  NOR2XL U1304 ( .A(N896), .B(n1792), .Y(psum3[2]) );
  NOR2XL U1305 ( .A(N896), .B(n1791), .Y(psum3[3]) );
  NOR2XL U1306 ( .A(N896), .B(n1790), .Y(psum3[4]) );
  NOR2XL U1307 ( .A(N896), .B(n1789), .Y(psum3[5]) );
  NOR2XL U1308 ( .A(N896), .B(n1788), .Y(psum3[6]) );
  NOR2XL U1309 ( .A(N892), .B(n1769), .Y(psum1[1]) );
  NOR2XL U1310 ( .A(N892), .B(n1768), .Y(psum1[2]) );
  NOR2XL U1311 ( .A(N892), .B(n1767), .Y(psum1[3]) );
  NOR2XL U1312 ( .A(N892), .B(n1766), .Y(psum1[4]) );
  NOR2XL U1313 ( .A(N892), .B(n1765), .Y(psum1[5]) );
  NOR2XL U1314 ( .A(N892), .B(n1764), .Y(psum1[6]) );
  NOR2XL U1315 ( .A(N894), .B(n1785), .Y(psum2[1]) );
  AO22X1 U1316 ( .A0(n1619), .A1(n1695), .B0(N261), .B1(n1620), .Y(n1502) );
  AO22X1 U1317 ( .A0(n1694), .A1(n1619), .B0(N260), .B1(n1620), .Y(n1503) );
  AO22X1 U1318 ( .A0(n1619), .A1(n1688), .B0(N269), .B1(n1620), .Y(n1493) );
  AO22X1 U1319 ( .A0(n1687), .A1(n1619), .B0(N268), .B1(n1620), .Y(n1494) );
  NOR2XL U1320 ( .A(N894), .B(n1779), .Y(psum2[7]) );
  NOR2XL U1321 ( .A(N896), .B(n1787), .Y(psum3[7]) );
  NOR2XL U1322 ( .A(N892), .B(n1763), .Y(psum1[7]) );
  NOR2XL U1323 ( .A(N898), .B(n1802), .Y(psum4[0]) );
  NOR2XL U1324 ( .A(N898), .B(n1801), .Y(psum4[1]) );
  NOR2XL U1325 ( .A(N898), .B(n1800), .Y(psum4[2]) );
  NOR2XL U1326 ( .A(N898), .B(n1799), .Y(psum4[3]) );
  NOR2XL U1327 ( .A(N898), .B(n1798), .Y(psum4[4]) );
  NOR2XL U1328 ( .A(N898), .B(n1797), .Y(psum4[5]) );
  NOR2XL U1329 ( .A(N898), .B(n1796), .Y(psum4[6]) );
  NOR2XL U1330 ( .A(N898), .B(n1795), .Y(psum4[7]) );
  CLKINVX1 U1331 ( .A(n1630), .Y(n1743) );
  AND2X2 U1332 ( .A(n1266), .B(n1267), .Y(n918) );
  NOR3X1 U1333 ( .A(n1624), .B(n1622), .C(n1623), .Y(n1267) );
  NOR3X1 U1334 ( .A(n1621), .B(n1625), .C(n1626), .Y(n1266) );
  NOR2BX1 U1335 ( .AN(n1198), .B(n1686), .Y(n1268) );
  NOR2BX1 U1336 ( .AN(n1014), .B(n1693), .Y(n1146) );
  NOR2X1 U1337 ( .A(n1628), .B(n1630), .Y(n1164) );
  NOR2X1 U1338 ( .A(n1629), .B(n1631), .Y(n1165) );
  NAND3X2 U1339 ( .A(n1628), .B(n1630), .C(n1197), .Y(n974) );
  NOR3BX1 U1340 ( .AN(n1272), .B(n785), .C(n1687), .Y(n1198) );
  NOR3BX1 U1341 ( .AN(n788), .B(n785), .C(n1694), .Y(n1014) );
  CLKINVX1 U1342 ( .A(n920), .Y(n1755) );
  CLKINVX1 U1343 ( .A(n923), .Y(n1756) );
  CLKINVX1 U1344 ( .A(n926), .Y(n1757) );
  CLKINVX1 U1345 ( .A(n929), .Y(n1758) );
  CLKINVX1 U1346 ( .A(n932), .Y(n1759) );
  CLKINVX1 U1347 ( .A(n935), .Y(n1760) );
  CLKINVX1 U1348 ( .A(n938), .Y(n1761) );
  CLKINVX1 U1349 ( .A(n954), .Y(n1762) );
  INVX3 U1350 ( .A(n941), .Y(n1906) );
  NAND3X1 U1351 ( .A(n1628), .B(n1630), .C(n1165), .Y(n970) );
  NAND2X1 U1352 ( .A(n1197), .B(n1164), .Y(n975) );
  INVX3 U1353 ( .A(n785), .Y(n1907) );
  NOR2X1 U1354 ( .A(index_a[2]), .B(n1691), .Y(n1153) );
  NOR2X1 U1355 ( .A(n1685), .B(n1683), .Y(n1275) );
  CLKINVX1 U1356 ( .A(n879), .Y(n1771) );
  CLKINVX1 U1357 ( .A(n882), .Y(n1772) );
  CLKINVX1 U1358 ( .A(n885), .Y(n1773) );
  CLKINVX1 U1359 ( .A(n888), .Y(n1774) );
  CLKINVX1 U1360 ( .A(n891), .Y(n1775) );
  CLKINVX1 U1361 ( .A(n894), .Y(n1776) );
  CLKINVX1 U1362 ( .A(n897), .Y(n1777) );
  CLKINVX1 U1363 ( .A(n900), .Y(n1778) );
  CLKBUFX3 U1364 ( .A(n1254), .Y(n1594) );
  NAND3X1 U1365 ( .A(n1682), .B(n1684), .C(n1268), .Y(n1254) );
  CLKBUFX3 U1366 ( .A(n840), .Y(n1678) );
  CLKBUFX3 U1367 ( .A(n840), .Y(n1679) );
  CLKBUFX3 U1368 ( .A(n841), .Y(n1676) );
  CLKBUFX3 U1369 ( .A(n844), .Y(n1672) );
  CLKBUFX3 U1370 ( .A(n1138), .Y(n1596) );
  NAND3BX1 U1371 ( .AN(n1627), .B(n918), .C(n1906), .Y(n1138) );
  INVX3 U1372 ( .A(n1692), .Y(n1691) );
  INVX3 U1373 ( .A(n1655), .Y(n1657) );
  AND2X2 U1374 ( .A(n1225), .B(n1197), .Y(n1571) );
  NAND2X1 U1375 ( .A(n1225), .B(n1165), .Y(n971) );
  NAND3X1 U1376 ( .A(n1629), .B(n1631), .C(n1164), .Y(n965) );
  CLKBUFX3 U1377 ( .A(n967), .Y(n1661) );
  NAND3X1 U1378 ( .A(n1629), .B(n1631), .C(n1225), .Y(n967) );
  CLKBUFX3 U1379 ( .A(n843), .Y(n1675) );
  CLKBUFX3 U1380 ( .A(n843), .Y(n1674) );
  CLKBUFX3 U1381 ( .A(n781), .Y(n1619) );
  NOR2X1 U1382 ( .A(n1509), .B(n1907), .Y(n781) );
  CLKBUFX3 U1383 ( .A(n844), .Y(n1673) );
  CLKBUFX3 U1384 ( .A(n841), .Y(n1677) );
  INVX3 U1385 ( .A(n1669), .Y(n1671) );
  INVX3 U1386 ( .A(n968), .Y(n1660) );
  OAI221XL U1387 ( .A0(n1762), .A1(n794), .B0(n795), .B1(n724), .C0(n796), .Y(
        n1283) );
  NAND2X1 U1388 ( .A(data_in_o[0]), .B(n797), .Y(n796) );
  OAI221XL U1389 ( .A0(n1761), .A1(n794), .B0(n795), .B1(n723), .C0(n798), .Y(
        n1284) );
  NAND2X1 U1390 ( .A(data_in_o[1]), .B(n797), .Y(n798) );
  OAI221XL U1391 ( .A0(n1760), .A1(n794), .B0(n795), .B1(n722), .C0(n799), .Y(
        n1285) );
  NAND2X1 U1392 ( .A(data_in_o[2]), .B(n1540), .Y(n799) );
  OAI221XL U1393 ( .A0(n1759), .A1(n794), .B0(n795), .B1(n721), .C0(n800), .Y(
        n1286) );
  NAND2X1 U1394 ( .A(data_in_o[3]), .B(n1540), .Y(n800) );
  OAI221XL U1395 ( .A0(n1758), .A1(n794), .B0(n795), .B1(n720), .C0(n801), .Y(
        n1287) );
  NAND2X1 U1396 ( .A(data_in_o[4]), .B(n797), .Y(n801) );
  OAI221XL U1397 ( .A0(n1757), .A1(n794), .B0(n795), .B1(n719), .C0(n802), .Y(
        n1288) );
  NAND2X1 U1398 ( .A(data_in_o[5]), .B(n1540), .Y(n802) );
  OAI221XL U1399 ( .A0(n1756), .A1(n794), .B0(n795), .B1(n718), .C0(n803), .Y(
        n1289) );
  NAND2X1 U1400 ( .A(data_in_o[6]), .B(n797), .Y(n803) );
  OAI221XL U1401 ( .A0(n1755), .A1(n794), .B0(n795), .B1(n717), .C0(n804), .Y(
        n1290) );
  NAND2X1 U1402 ( .A(data_in_o[7]), .B(n1540), .Y(n804) );
  NAND2X1 U1403 ( .A(data_in_o[8]), .B(n1540), .Y(n811) );
  NAND2X1 U1404 ( .A(data_in_o[9]), .B(n1540), .Y(n812) );
  NAND2X1 U1405 ( .A(data_in_o[10]), .B(n1540), .Y(n813) );
  NAND2X1 U1406 ( .A(data_in_o[11]), .B(n1540), .Y(n814) );
  NAND2X1 U1407 ( .A(data_in_o[12]), .B(n1540), .Y(n815) );
  NAND2X1 U1408 ( .A(data_in_o[13]), .B(n1540), .Y(n816) );
  NAND2X1 U1409 ( .A(data_in_o[14]), .B(n1540), .Y(n817) );
  NAND2X1 U1410 ( .A(data_in_o[15]), .B(n797), .Y(n818) );
  OAI2BB2XL U1411 ( .B0(n1631), .B1(n1572), .A0N(n1743), .A1N(N780), .Y(n1707)
         );
  XNOR2X1 U1412 ( .A(n[0]), .B(N785), .Y(n1572) );
  OAI2BB2XL U1413 ( .B0(n839), .B1(n1618), .A0N(data_in_o[24]), .A1N(n797), 
        .Y(n1299) );
  AOI221XL U1414 ( .A0(w42[0]), .A1(n1679), .B0(w41[0]), .B1(n1677), .C0(n842), 
        .Y(n839) );
  OAI2BB2XL U1415 ( .B0(n1802), .B1(n1674), .A0N(w43[0]), .A1N(n1673), .Y(n842) );
  OAI2BB2XL U1416 ( .B0(n845), .B1(n1618), .A0N(data_in_o[25]), .A1N(n797), 
        .Y(n1300) );
  AOI221XL U1417 ( .A0(w42[1]), .A1(n1679), .B0(w41[1]), .B1(n1677), .C0(n846), 
        .Y(n845) );
  OAI2BB2XL U1418 ( .B0(n1801), .B1(n1674), .A0N(w43[1]), .A1N(n1673), .Y(n846) );
  OAI2BB2XL U1419 ( .B0(n847), .B1(n1618), .A0N(data_in_o[26]), .A1N(n797), 
        .Y(n1301) );
  AOI221XL U1420 ( .A0(w42[2]), .A1(n1679), .B0(w41[2]), .B1(n1677), .C0(n848), 
        .Y(n847) );
  OAI2BB2XL U1421 ( .B0(n1800), .B1(n1674), .A0N(w43[2]), .A1N(n1672), .Y(n848) );
  OAI2BB2XL U1422 ( .B0(n849), .B1(n1618), .A0N(data_in_o[27]), .A1N(n797), 
        .Y(n1302) );
  AOI221XL U1423 ( .A0(w42[3]), .A1(n1679), .B0(w41[3]), .B1(n1677), .C0(n850), 
        .Y(n849) );
  OAI2BB2XL U1424 ( .B0(n1799), .B1(n1674), .A0N(w43[3]), .A1N(n1673), .Y(n850) );
  OAI2BB2XL U1425 ( .B0(n851), .B1(n1618), .A0N(data_in_o[28]), .A1N(n797), 
        .Y(n1303) );
  AOI221XL U1426 ( .A0(w42[4]), .A1(n1678), .B0(w41[4]), .B1(n1677), .C0(n852), 
        .Y(n851) );
  OAI2BB2XL U1427 ( .B0(n1798), .B1(n1674), .A0N(w43[4]), .A1N(n1672), .Y(n852) );
  OAI2BB2XL U1428 ( .B0(n853), .B1(n1618), .A0N(data_in_o[29]), .A1N(n797), 
        .Y(n1304) );
  AOI221XL U1429 ( .A0(w42[5]), .A1(n1679), .B0(w41[5]), .B1(n1677), .C0(n854), 
        .Y(n853) );
  OAI2BB2XL U1430 ( .B0(n1797), .B1(n1674), .A0N(w43[5]), .A1N(n1673), .Y(n854) );
  OAI2BB2XL U1431 ( .B0(n855), .B1(n1618), .A0N(data_in_o[30]), .A1N(n797), 
        .Y(n1305) );
  AOI221XL U1432 ( .A0(w42[6]), .A1(n1679), .B0(w41[6]), .B1(n1677), .C0(n856), 
        .Y(n855) );
  OAI2BB2XL U1433 ( .B0(n1796), .B1(n1674), .A0N(w43[6]), .A1N(n1673), .Y(n856) );
  OAI2BB2XL U1434 ( .B0(n857), .B1(n1618), .A0N(data_in_o[31]), .A1N(n797), 
        .Y(n1306) );
  AOI221XL U1435 ( .A0(w42[7]), .A1(n1679), .B0(w41[7]), .B1(n1677), .C0(n858), 
        .Y(n857) );
  OAI2BB2XL U1436 ( .B0(n1795), .B1(n1674), .A0N(w43[7]), .A1N(n1673), .Y(n858) );
  CLKINVX1 U1437 ( .A(n828), .Y(n1749) );
  CLKINVX1 U1438 ( .A(n834), .Y(n1750) );
  CLKINVX1 U1439 ( .A(n836), .Y(n1751) );
  OAI222XL U1440 ( .A0(n903), .A1(n733), .B0(n1755), .B1(n904), .C0(n1617), 
        .C1(n717), .Y(n1315) );
  OAI222XL U1441 ( .A0(n903), .A1(n734), .B0(n1756), .B1(n904), .C0(n1617), 
        .C1(n718), .Y(n1316) );
  OAI222XL U1442 ( .A0(n903), .A1(n735), .B0(n1757), .B1(n904), .C0(n1617), 
        .C1(n719), .Y(n1317) );
  OAI222XL U1443 ( .A0(n903), .A1(n736), .B0(n1758), .B1(n904), .C0(n1617), 
        .C1(n720), .Y(n1318) );
  OAI222XL U1444 ( .A0(n903), .A1(n737), .B0(n1759), .B1(n904), .C0(n1617), 
        .C1(n721), .Y(n1319) );
  OAI222XL U1445 ( .A0(n903), .A1(n738), .B0(n1760), .B1(n904), .C0(n1617), 
        .C1(n722), .Y(n1320) );
  OAI222XL U1446 ( .A0(n903), .A1(n739), .B0(n1761), .B1(n904), .C0(n1617), 
        .C1(n723), .Y(n1321) );
  OAI222XL U1447 ( .A0(n903), .A1(n740), .B0(n1762), .B1(n904), .C0(n1617), 
        .C1(n724), .Y(n1322) );
  OAI222XL U1448 ( .A0(n1615), .A1(n725), .B0(n1771), .B1(n1616), .C0(n1614), 
        .C1(n709), .Y(n1307) );
  OAI222XL U1449 ( .A0(n1615), .A1(n726), .B0(n1772), .B1(n1616), .C0(n1542), 
        .C1(n710), .Y(n1308) );
  OAI222XL U1450 ( .A0(n1615), .A1(n727), .B0(n1773), .B1(n1616), .C0(n1542), 
        .C1(n711), .Y(n1309) );
  OAI222XL U1451 ( .A0(n1615), .A1(n728), .B0(n1774), .B1(n1616), .C0(n1542), 
        .C1(n712), .Y(n1310) );
  OAI222XL U1452 ( .A0(n1615), .A1(n729), .B0(n1775), .B1(n1616), .C0(n1542), 
        .C1(n713), .Y(n1311) );
  OAI222XL U1453 ( .A0(n1615), .A1(n730), .B0(n1776), .B1(n1616), .C0(n1542), 
        .C1(n714), .Y(n1312) );
  OAI222XL U1454 ( .A0(n1615), .A1(n731), .B0(n1777), .B1(n1616), .C0(n1542), 
        .C1(n715), .Y(n1313) );
  OAI222XL U1455 ( .A0(n1615), .A1(n732), .B0(n1778), .B1(n1616), .C0(n1542), 
        .C1(n716), .Y(n1314) );
  OAI222XL U1456 ( .A0(n1615), .A1(n701), .B0(n1755), .B1(n1616), .C0(n1542), 
        .C1(n733), .Y(n1323) );
  OAI222XL U1457 ( .A0(n1615), .A1(n702), .B0(n1756), .B1(n1616), .C0(n1542), 
        .C1(n734), .Y(n1324) );
  OAI222XL U1458 ( .A0(n1615), .A1(n707), .B0(n1761), .B1(n877), .C0(n1542), 
        .C1(n739), .Y(n1329) );
  XOR2X1 U1459 ( .A(n[3]), .B(\add_357_2/carry[4] ), .Y(N789) );
  OAI2BB2XL U1460 ( .B0(n1631), .B1(N785), .A0N(n1743), .A1N(N712), .Y(n1718)
         );
  AND2X2 U1461 ( .A(n[3]), .B(\add_357_2/carry[4] ), .Y(n1573) );
  NAND4X1 U1462 ( .A(n948), .B(n918), .C(n949), .D(n950), .Y(n909) );
  XOR2X1 U1463 ( .A(n700), .B(N785), .Y(n948) );
  XNOR2X1 U1464 ( .A(n1627), .B(n1576), .Y(n949) );
  NOR3X1 U1465 ( .A(n951), .B(n952), .C(n953), .Y(n950) );
  XOR2X1 U1466 ( .A(n700), .B(n1529), .Y(n942) );
  XNOR2X1 U1467 ( .A(n1627), .B(N722), .Y(n943) );
  XOR2X1 U1468 ( .A(n1628), .B(N727), .Y(n951) );
  XOR2X1 U1469 ( .A(n1629), .B(N726), .Y(n952) );
  XNOR2X1 U1470 ( .A(n1628), .B(N733), .Y(n916) );
  XNOR2X1 U1471 ( .A(n1629), .B(N732), .Y(n914) );
  XOR2X1 U1472 ( .A(n699), .B(N731), .Y(n917) );
  XOR2X1 U1473 ( .A(n1627), .B(n1577), .Y(n919) );
  OAI21XL U1474 ( .A0(n1855), .A1(n1278), .B0(n1279), .Y(N252) );
  AO22X1 U1475 ( .A0(N244), .A1(n1276), .B0(n1854), .B1(n1277), .Y(N254) );
  CLKINVX1 U1476 ( .A(\sub_142/carry[4] ), .Y(N244) );
  CLKBUFX3 U1477 ( .A(counter[4]), .Y(n1627) );
  CLKBUFX3 U1478 ( .A(counter[1]), .Y(n1630) );
  CLKBUFX3 U1479 ( .A(counter[0]), .Y(n1631) );
  CLKBUFX3 U1480 ( .A(counter[5]), .Y(n1626) );
  CLKBUFX3 U1481 ( .A(counter[6]), .Y(n1625) );
  CLKBUFX3 U1482 ( .A(counter[7]), .Y(n1624) );
  CLKBUFX3 U1483 ( .A(counter[9]), .Y(n1622) );
  AO22X1 U1484 ( .A0(n1619), .A1(index_b[7]), .B0(N272), .B1(n1620), .Y(n1498)
         );
  AO22X1 U1485 ( .A0(n1619), .A1(index_a[7]), .B0(N264), .B1(n1620), .Y(n1508)
         );
  CLKBUFX3 U1486 ( .A(counter[8]), .Y(n1623) );
  AO22X1 U1487 ( .A0(N243), .A1(n1276), .B0(n1854), .B1(n1277), .Y(N253) );
  AO22X1 U1488 ( .A0(n1619), .A1(index_a[6]), .B0(N263), .B1(n1620), .Y(n1500)
         );
  AO22X1 U1489 ( .A0(n1619), .A1(index_a[5]), .B0(N262), .B1(n1620), .Y(n1501)
         );
  AO22X1 U1490 ( .A0(n1619), .A1(index_b[6]), .B0(N271), .B1(n1620), .Y(n1491)
         );
  AO22X1 U1491 ( .A0(n1619), .A1(index_b[5]), .B0(N270), .B1(n1620), .Y(n1492)
         );
  CLKBUFX3 U1492 ( .A(counter[10]), .Y(n1621) );
  OAI221XL U1493 ( .A0(load_en), .A1(n225), .B0(n163), .B1(n741), .C0(n779), 
        .Y(next_state[0]) );
  AOI21X1 U1494 ( .A0(start), .A1(n1509), .B0(N912), .Y(n779) );
  NOR2X1 U1495 ( .A(n163), .B(n225), .Y(N912) );
  OAI2BB2XL U1496 ( .B0(n785), .B1(n786), .A0N(load_en), .A1N(n1619), .Y(n1507) );
  OAI222XL U1497 ( .A0(n1670), .A1(n361), .B0(n1666), .B1(n369), .C0(n1665), 
        .C1(n257), .Y(n1012) );
  OAI222XL U1498 ( .A0(n1670), .A1(n360), .B0(n1666), .B1(n368), .C0(n1665), 
        .C1(n256), .Y(n1005) );
  OAI222XL U1499 ( .A0(n1670), .A1(n359), .B0(n1667), .B1(n367), .C0(n1665), 
        .C1(n255), .Y(n1000) );
  OAI222XL U1500 ( .A0(n1669), .A1(n358), .B0(n1667), .B1(n366), .C0(n1665), 
        .C1(n254), .Y(n995) );
  OAI222XL U1501 ( .A0(n1670), .A1(n357), .B0(n1667), .B1(n365), .C0(n1665), 
        .C1(n253), .Y(n990) );
  OAI222XL U1502 ( .A0(n1670), .A1(n356), .B0(n1667), .B1(n364), .C0(n1665), 
        .C1(n252), .Y(n985) );
  OAI222XL U1503 ( .A0(n1670), .A1(n355), .B0(n1667), .B1(n363), .C0(n1665), 
        .C1(n251), .Y(n980) );
  OAI222XL U1504 ( .A0(n1670), .A1(n354), .B0(n1667), .B1(n362), .C0(n1665), 
        .C1(n250), .Y(n963) );
  OAI222XL U1505 ( .A0(n1662), .A1(n385), .B0(n1658), .B1(n489), .C0(n969), 
        .C1(n377), .Y(n1011) );
  OAI222XL U1506 ( .A0(n1662), .A1(n384), .B0(n1658), .B1(n488), .C0(n969), 
        .C1(n376), .Y(n1004) );
  OAI222XL U1507 ( .A0(n1662), .A1(n383), .B0(n1658), .B1(n487), .C0(n969), 
        .C1(n375), .Y(n999) );
  OAI222XL U1508 ( .A0(n1661), .A1(n382), .B0(n1658), .B1(n486), .C0(n1655), 
        .C1(n374), .Y(n994) );
  OAI222XL U1509 ( .A0(n1595), .A1(n501), .B0(n1652), .B1(n245), .C0(n1649), 
        .C1(n493), .Y(n988) );
  OAI222XL U1510 ( .A0(n1595), .A1(n500), .B0(n1652), .B1(n244), .C0(n1649), 
        .C1(n492), .Y(n983) );
  OAI222XL U1511 ( .A0(n1595), .A1(n499), .B0(n1652), .B1(n243), .C0(n1649), 
        .C1(n491), .Y(n978) );
  OAI222XL U1512 ( .A0(n1595), .A1(n498), .B0(n1652), .B1(n242), .C0(n1649), 
        .C1(n490), .Y(n961) );
  OAI211X1 U1513 ( .A0(n1779), .A1(n1675), .B0(n880), .C0(n881), .Y(n879) );
  NAND2X1 U1514 ( .A(w23[7]), .B(n1673), .Y(n880) );
  AOI22X1 U1515 ( .A0(w22[7]), .A1(n1679), .B0(w21[7]), .B1(n1677), .Y(n881)
         );
  OAI211X1 U1516 ( .A0(n1780), .A1(n1675), .B0(n883), .C0(n884), .Y(n882) );
  NAND2X1 U1517 ( .A(w23[6]), .B(n1673), .Y(n883) );
  AOI22X1 U1518 ( .A0(w22[6]), .A1(n1679), .B0(w21[6]), .B1(n1677), .Y(n884)
         );
  OAI211X1 U1519 ( .A0(n1781), .A1(n1675), .B0(n886), .C0(n887), .Y(n885) );
  NAND2X1 U1520 ( .A(w23[5]), .B(n1673), .Y(n886) );
  AOI22X1 U1521 ( .A0(w22[5]), .A1(n1679), .B0(w21[5]), .B1(n1677), .Y(n887)
         );
  OAI211X1 U1522 ( .A0(n1782), .A1(n1675), .B0(n889), .C0(n890), .Y(n888) );
  NAND2X1 U1523 ( .A(w23[4]), .B(n1673), .Y(n889) );
  AOI22X1 U1524 ( .A0(w22[4]), .A1(n1678), .B0(w21[4]), .B1(n1677), .Y(n890)
         );
  OAI211X1 U1525 ( .A0(n1783), .A1(n1675), .B0(n892), .C0(n893), .Y(n891) );
  NAND2X1 U1526 ( .A(w23[3]), .B(n1672), .Y(n892) );
  AOI22X1 U1527 ( .A0(w22[3]), .A1(n1678), .B0(w21[3]), .B1(n1676), .Y(n893)
         );
  OAI211X1 U1528 ( .A0(n1784), .A1(n1675), .B0(n895), .C0(n896), .Y(n894) );
  NAND2X1 U1529 ( .A(w23[2]), .B(n1672), .Y(n895) );
  AOI22X1 U1530 ( .A0(w22[2]), .A1(n1678), .B0(w21[2]), .B1(n1676), .Y(n896)
         );
  OAI211X1 U1531 ( .A0(n1785), .A1(n1675), .B0(n898), .C0(n899), .Y(n897) );
  NAND2X1 U1532 ( .A(w23[1]), .B(n1672), .Y(n898) );
  AOI22X1 U1533 ( .A0(w22[1]), .A1(n1678), .B0(w21[1]), .B1(n1676), .Y(n899)
         );
  OAI211X1 U1534 ( .A0(n1763), .A1(n1675), .B0(n921), .C0(n922), .Y(n920) );
  NAND2X1 U1535 ( .A(w13[7]), .B(n1672), .Y(n921) );
  AOI22X1 U1536 ( .A0(w12[7]), .A1(n1678), .B0(w11[7]), .B1(n1676), .Y(n922)
         );
  OAI211X1 U1537 ( .A0(n1764), .A1(n1675), .B0(n924), .C0(n925), .Y(n923) );
  NAND2X1 U1538 ( .A(w13[6]), .B(n1672), .Y(n924) );
  AOI22X1 U1539 ( .A0(w12[6]), .A1(n1678), .B0(w11[6]), .B1(n1676), .Y(n925)
         );
  OAI211X1 U1540 ( .A0(n1765), .A1(n1675), .B0(n927), .C0(n928), .Y(n926) );
  NAND2X1 U1541 ( .A(w13[5]), .B(n1672), .Y(n927) );
  AOI22X1 U1542 ( .A0(w12[5]), .A1(n1678), .B0(w11[5]), .B1(n1676), .Y(n928)
         );
  OAI211X1 U1543 ( .A0(n1766), .A1(n1675), .B0(n930), .C0(n931), .Y(n929) );
  NAND2X1 U1544 ( .A(w13[4]), .B(n1672), .Y(n930) );
  AOI22X1 U1545 ( .A0(w12[4]), .A1(n1678), .B0(w11[4]), .B1(n1676), .Y(n931)
         );
  OAI211X1 U1546 ( .A0(n1767), .A1(n1675), .B0(n933), .C0(n934), .Y(n932) );
  NAND2X1 U1547 ( .A(w13[3]), .B(n1672), .Y(n933) );
  AOI22X1 U1548 ( .A0(w12[3]), .A1(n1678), .B0(w11[3]), .B1(n1676), .Y(n934)
         );
  OAI211X1 U1549 ( .A0(n1768), .A1(n1675), .B0(n936), .C0(n937), .Y(n935) );
  NAND2X1 U1550 ( .A(w13[2]), .B(n1672), .Y(n936) );
  AOI22X1 U1551 ( .A0(w12[2]), .A1(n1678), .B0(w11[2]), .B1(n1676), .Y(n937)
         );
  OAI211X1 U1552 ( .A0(n1769), .A1(n1675), .B0(n939), .C0(n940), .Y(n938) );
  NAND2X1 U1553 ( .A(w13[1]), .B(n1672), .Y(n939) );
  AOI22X1 U1554 ( .A0(w12[1]), .A1(n1678), .B0(w11[1]), .B1(n1676), .Y(n940)
         );
  OAI211X1 U1555 ( .A0(n1787), .A1(n1674), .B0(n860), .C0(n861), .Y(n837) );
  NAND2X1 U1556 ( .A(w33[7]), .B(n1673), .Y(n860) );
  AOI22X1 U1557 ( .A0(w32[7]), .A1(n1679), .B0(w31[7]), .B1(n1676), .Y(n861)
         );
  OAI211X1 U1558 ( .A0(n1788), .A1(n1674), .B0(n862), .C0(n863), .Y(n835) );
  NAND2X1 U1559 ( .A(w33[6]), .B(n1673), .Y(n862) );
  AOI22X1 U1560 ( .A0(w32[6]), .A1(n1679), .B0(w31[6]), .B1(n1677), .Y(n863)
         );
  OAI211X1 U1561 ( .A0(n1789), .A1(n1674), .B0(n864), .C0(n865), .Y(n833) );
  NAND2X1 U1562 ( .A(w33[5]), .B(n1673), .Y(n864) );
  AOI22X1 U1563 ( .A0(w32[5]), .A1(n1679), .B0(w31[5]), .B1(n1677), .Y(n865)
         );
  OAI211X1 U1564 ( .A0(n1790), .A1(n1674), .B0(n866), .C0(n867), .Y(n831) );
  NAND2X1 U1565 ( .A(w33[4]), .B(n1673), .Y(n866) );
  AOI22X1 U1566 ( .A0(w32[4]), .A1(n1679), .B0(w31[4]), .B1(n1677), .Y(n867)
         );
  OAI211X1 U1567 ( .A0(n1791), .A1(n1674), .B0(n868), .C0(n869), .Y(n829) );
  NAND2X1 U1568 ( .A(w33[3]), .B(n1673), .Y(n868) );
  AOI22X1 U1569 ( .A0(w32[3]), .A1(n1679), .B0(w31[3]), .B1(n1676), .Y(n869)
         );
  NAND2X1 U1570 ( .A(w33[2]), .B(n1673), .Y(n870) );
  AOI22X1 U1571 ( .A0(w32[2]), .A1(n1679), .B0(w31[2]), .B1(n1677), .Y(n871)
         );
  OAI211X1 U1572 ( .A0(n1793), .A1(n1675), .B0(n872), .C0(n873), .Y(n825) );
  NAND2X1 U1573 ( .A(w33[1]), .B(n1673), .Y(n872) );
  AOI22X1 U1574 ( .A0(w32[1]), .A1(n1679), .B0(w31[1]), .B1(n1677), .Y(n873)
         );
  OAI211X1 U1575 ( .A0(n1794), .A1(n1675), .B0(n874), .C0(n875), .Y(n823) );
  NAND2X1 U1576 ( .A(w33[0]), .B(n1673), .Y(n874) );
  AOI22X1 U1577 ( .A0(w32[0]), .A1(n1679), .B0(w31[0]), .B1(n1677), .Y(n875)
         );
  OAI222XL U1578 ( .A0(n1599), .A1(n553), .B0(n1600), .B1(n593), .C0(n1598), 
        .C1(n666), .Y(n1466) );
  OAI222XL U1579 ( .A0(n1599), .A1(n552), .B0(n1600), .B1(n592), .C0(n1598), 
        .C1(n665), .Y(n1465) );
  OAI222XL U1580 ( .A0(n1599), .A1(n551), .B0(n1600), .B1(n591), .C0(n1598), 
        .C1(n664), .Y(n1464) );
  OAI222XL U1581 ( .A0(n1599), .A1(n550), .B0(n1600), .B1(n590), .C0(n1598), 
        .C1(n663), .Y(n1463) );
  OAI222XL U1582 ( .A0(n1599), .A1(n549), .B0(n1600), .B1(n589), .C0(n1598), 
        .C1(n662), .Y(n1462) );
  OAI222XL U1583 ( .A0(n1599), .A1(n548), .B0(n1600), .B1(n588), .C0(n1598), 
        .C1(n661), .Y(n1461) );
  OAI222XL U1584 ( .A0(n1599), .A1(n547), .B0(n1600), .B1(n587), .C0(n1598), 
        .C1(n660), .Y(n1460) );
  OAI222XL U1585 ( .A0(n1599), .A1(n546), .B0(n1600), .B1(n586), .C0(n1598), 
        .C1(n659), .Y(n1459) );
  OAI222XL U1586 ( .A0(n1602), .A1(n585), .B0(n1603), .B1(n529), .C0(n1601), 
        .C1(n650), .Y(n1442) );
  OAI222XL U1587 ( .A0(n1602), .A1(n584), .B0(n1603), .B1(n528), .C0(n1601), 
        .C1(n649), .Y(n1441) );
  OAI222XL U1588 ( .A0(n1602), .A1(n583), .B0(n1603), .B1(n527), .C0(n1601), 
        .C1(n648), .Y(n1440) );
  OAI222XL U1589 ( .A0(n1602), .A1(n582), .B0(n1603), .B1(n526), .C0(n1601), 
        .C1(n647), .Y(n1439) );
  OAI222XL U1590 ( .A0(n1602), .A1(n581), .B0(n1603), .B1(n525), .C0(n1601), 
        .C1(n646), .Y(n1438) );
  OAI222XL U1591 ( .A0(n1602), .A1(n580), .B0(n1603), .B1(n524), .C0(n1601), 
        .C1(n645), .Y(n1437) );
  OAI222XL U1592 ( .A0(n1602), .A1(n579), .B0(n1603), .B1(n523), .C0(n1601), 
        .C1(n644), .Y(n1436) );
  OAI222XL U1593 ( .A0(n1602), .A1(n578), .B0(n1603), .B1(n522), .C0(n1601), 
        .C1(n643), .Y(n1435) );
  OAI222XL U1594 ( .A0(n1602), .A1(n577), .B0(n1603), .B1(n537), .C0(n1601), 
        .C1(n658), .Y(n1450) );
  OAI222XL U1595 ( .A0(n1602), .A1(n576), .B0(n1603), .B1(n536), .C0(n1601), 
        .C1(n657), .Y(n1449) );
  OAI222XL U1596 ( .A0(n1602), .A1(n575), .B0(n1603), .B1(n535), .C0(n1601), 
        .C1(n656), .Y(n1448) );
  OAI222XL U1597 ( .A0(n1602), .A1(n574), .B0(n1603), .B1(n534), .C0(n1601), 
        .C1(n655), .Y(n1447) );
  OAI222XL U1598 ( .A0(n1602), .A1(n573), .B0(n1603), .B1(n533), .C0(n1601), 
        .C1(n654), .Y(n1446) );
  OAI222XL U1599 ( .A0(n1602), .A1(n572), .B0(n1603), .B1(n532), .C0(n1601), 
        .C1(n653), .Y(n1445) );
  OAI222XL U1600 ( .A0(n1602), .A1(n571), .B0(n1603), .B1(n531), .C0(n1601), 
        .C1(n652), .Y(n1444) );
  OAI222XL U1601 ( .A0(n1602), .A1(n570), .B0(n1603), .B1(n530), .C0(n1601), 
        .C1(n651), .Y(n1443) );
  OAI222XL U1602 ( .A0(n1199), .A1(n569), .B0(n1200), .B1(n521), .C0(n1605), 
        .C1(n642), .Y(n1434) );
  OAI222XL U1603 ( .A0(n1199), .A1(n568), .B0(n1200), .B1(n520), .C0(n1605), 
        .C1(n641), .Y(n1433) );
  OAI222XL U1604 ( .A0(n1199), .A1(n567), .B0(n1200), .B1(n519), .C0(n1605), 
        .C1(n640), .Y(n1432) );
  OAI222XL U1605 ( .A0(n1199), .A1(n566), .B0(n1200), .B1(n518), .C0(n1605), 
        .C1(n639), .Y(n1431) );
  OAI222XL U1606 ( .A0(n1199), .A1(n565), .B0(n1200), .B1(n517), .C0(n1605), 
        .C1(n638), .Y(n1430) );
  OAI222XL U1607 ( .A0(n1199), .A1(n564), .B0(n1200), .B1(n516), .C0(n1605), 
        .C1(n637), .Y(n1429) );
  OAI222XL U1608 ( .A0(n1199), .A1(n563), .B0(n1200), .B1(n515), .C0(n1605), 
        .C1(n636), .Y(n1428) );
  OAI222XL U1609 ( .A0(n1199), .A1(n562), .B0(n1200), .B1(n514), .C0(n1605), 
        .C1(n635), .Y(n1427) );
  OAI222XL U1610 ( .A0(n1263), .A1(n561), .B0(n1264), .B1(n609), .C0(n1597), 
        .C1(n682), .Y(n1482) );
  OAI222XL U1611 ( .A0(n1263), .A1(n560), .B0(n1264), .B1(n608), .C0(n1597), 
        .C1(n681), .Y(n1481) );
  OAI222XL U1612 ( .A0(n1263), .A1(n559), .B0(n1264), .B1(n607), .C0(n1597), 
        .C1(n680), .Y(n1480) );
  OAI222XL U1613 ( .A0(n1263), .A1(n558), .B0(n1264), .B1(n606), .C0(n1597), 
        .C1(n679), .Y(n1479) );
  OAI222XL U1614 ( .A0(n1263), .A1(n557), .B0(n1264), .B1(n605), .C0(n1597), 
        .C1(n678), .Y(n1478) );
  OAI222XL U1615 ( .A0(n1263), .A1(n556), .B0(n1264), .B1(n604), .C0(n1597), 
        .C1(n677), .Y(n1477) );
  OAI222XL U1616 ( .A0(n1263), .A1(n555), .B0(n1264), .B1(n603), .C0(n1597), 
        .C1(n676), .Y(n1476) );
  OAI222XL U1617 ( .A0(n1263), .A1(n554), .B0(n1264), .B1(n602), .C0(n1597), 
        .C1(n675), .Y(n1475) );
  OAI222XL U1618 ( .A0(n1599), .A1(n545), .B0(n1600), .B1(n601), .C0(n1598), 
        .C1(n674), .Y(n1458) );
  OAI222XL U1619 ( .A0(n1599), .A1(n544), .B0(n1600), .B1(n600), .C0(n1598), 
        .C1(n673), .Y(n1457) );
  OAI222XL U1620 ( .A0(n1599), .A1(n543), .B0(n1600), .B1(n599), .C0(n1598), 
        .C1(n672), .Y(n1456) );
  OAI222XL U1621 ( .A0(n1599), .A1(n542), .B0(n1600), .B1(n598), .C0(n1598), 
        .C1(n671), .Y(n1455) );
  OAI222XL U1622 ( .A0(n1599), .A1(n541), .B0(n1600), .B1(n597), .C0(n1598), 
        .C1(n670), .Y(n1454) );
  OAI222XL U1623 ( .A0(n1599), .A1(n540), .B0(n1600), .B1(n596), .C0(n1598), 
        .C1(n669), .Y(n1453) );
  OAI222XL U1624 ( .A0(n1599), .A1(n539), .B0(n1600), .B1(n595), .C0(n1598), 
        .C1(n668), .Y(n1452) );
  OAI222XL U1625 ( .A0(n1599), .A1(n538), .B0(n1600), .B1(n594), .C0(n1598), 
        .C1(n667), .Y(n1451) );
  NOR3X1 U1626 ( .A(l[5]), .B(l[4]), .C(l[3]), .Y(n957) );
  OAI22XL U1627 ( .A0(n1664), .A1(n305), .B0(n1670), .B1(n313), .Y(n1099) );
  OAI22XL U1628 ( .A0(n1664), .A1(n304), .B0(n1670), .B1(n312), .Y(n1094) );
  OAI22XL U1629 ( .A0(n1664), .A1(n303), .B0(n1670), .B1(n311), .Y(n1089) );
  OAI22XL U1630 ( .A0(n1664), .A1(n302), .B0(n1670), .B1(n310), .Y(n1084) );
  OAI22XL U1631 ( .A0(n1664), .A1(n301), .B0(n1670), .B1(n309), .Y(n1079) );
  OAI22XL U1632 ( .A0(n1665), .A1(n300), .B0(n1669), .B1(n308), .Y(n1074) );
  OAI22XL U1633 ( .A0(n1665), .A1(n299), .B0(n1669), .B1(n307), .Y(n1069) );
  OAI22XL U1634 ( .A0(n1665), .A1(n298), .B0(n1669), .B1(n306), .Y(n1064) );
  OAI22XL U1635 ( .A0(n1665), .A1(n281), .B0(n1669), .B1(n289), .Y(n1056) );
  OAI22XL U1636 ( .A0(n1665), .A1(n280), .B0(n964), .B1(n288), .Y(n1050) );
  OAI22XL U1637 ( .A0(n1665), .A1(n279), .B0(n964), .B1(n287), .Y(n1045) );
  OAI22XL U1638 ( .A0(n1665), .A1(n278), .B0(n964), .B1(n286), .Y(n1040) );
  OAI22XL U1639 ( .A0(n1665), .A1(n277), .B0(n964), .B1(n285), .Y(n1035) );
  OAI22XL U1640 ( .A0(n1665), .A1(n276), .B0(n964), .B1(n284), .Y(n1030) );
  OAI22XL U1641 ( .A0(n1665), .A1(n275), .B0(n964), .B1(n283), .Y(n1025) );
  OAI22XL U1642 ( .A0(n1665), .A1(n274), .B0(n1669), .B1(n282), .Y(n1020) );
  OAI22XL U1643 ( .A0(n1664), .A1(n329), .B0(n1670), .B1(n337), .Y(n1144) );
  OAI22XL U1644 ( .A0(n1664), .A1(n328), .B0(n1670), .B1(n336), .Y(n1136) );
  OAI22XL U1645 ( .A0(n1664), .A1(n327), .B0(n1670), .B1(n335), .Y(n1131) );
  OAI22XL U1646 ( .A0(n1664), .A1(n326), .B0(n1670), .B1(n334), .Y(n1126) );
  OAI22XL U1647 ( .A0(n1664), .A1(n325), .B0(n1670), .B1(n333), .Y(n1121) );
  OAI22XL U1648 ( .A0(n1664), .A1(n324), .B0(n1670), .B1(n332), .Y(n1116) );
  OAI22XL U1649 ( .A0(n1664), .A1(n323), .B0(n1670), .B1(n331), .Y(n1111) );
  OAI22XL U1650 ( .A0(n1664), .A1(n322), .B0(n1670), .B1(n330), .Y(n1106) );
  OAI22XL U1651 ( .A0(n1662), .A1(n433), .B0(n1658), .B1(n441), .Y(n1097) );
  OAI22XL U1652 ( .A0(n1662), .A1(n432), .B0(n1658), .B1(n440), .Y(n1092) );
  OAI22XL U1653 ( .A0(n1662), .A1(n431), .B0(n1658), .B1(n439), .Y(n1087) );
  OAI22XL U1654 ( .A0(n1662), .A1(n430), .B0(n1658), .B1(n438), .Y(n1082) );
  OAI22XL U1655 ( .A0(n1662), .A1(n429), .B0(n1658), .B1(n437), .Y(n1077) );
  OAI22XL U1656 ( .A0(n1661), .A1(n428), .B0(n1658), .B1(n436), .Y(n1072) );
  OAI22XL U1657 ( .A0(n1661), .A1(n427), .B0(n1658), .B1(n435), .Y(n1067) );
  OAI22XL U1658 ( .A0(n1661), .A1(n426), .B0(n1658), .B1(n434), .Y(n1062) );
  OAI22XL U1659 ( .A0(n1661), .A1(n409), .B0(n1658), .B1(n417), .Y(n1054) );
  OAI22XL U1660 ( .A0(n1661), .A1(n408), .B0(n1658), .B1(n416), .Y(n1048) );
  OAI22XL U1661 ( .A0(n1661), .A1(n407), .B0(n1658), .B1(n415), .Y(n1043) );
  OAI22XL U1662 ( .A0(n967), .A1(n406), .B0(n1658), .B1(n414), .Y(n1038) );
  OAI22XL U1663 ( .A0(n967), .A1(n405), .B0(n1658), .B1(n413), .Y(n1033) );
  OAI22XL U1664 ( .A0(n967), .A1(n404), .B0(n1658), .B1(n412), .Y(n1028) );
  OAI22XL U1665 ( .A0(n967), .A1(n403), .B0(n1658), .B1(n411), .Y(n1023) );
  OAI22XL U1666 ( .A0(n967), .A1(n402), .B0(n1658), .B1(n410), .Y(n1018) );
  OAI22XL U1667 ( .A0(n1662), .A1(n457), .B0(n1658), .B1(n465), .Y(n1142) );
  OAI22XL U1668 ( .A0(n1662), .A1(n456), .B0(n1659), .B1(n464), .Y(n1134) );
  OAI22XL U1669 ( .A0(n1662), .A1(n455), .B0(n1659), .B1(n463), .Y(n1129) );
  OAI22XL U1670 ( .A0(n1662), .A1(n454), .B0(n968), .B1(n462), .Y(n1124) );
  OAI22XL U1671 ( .A0(n1662), .A1(n453), .B0(n968), .B1(n461), .Y(n1119) );
  OAI22XL U1672 ( .A0(n1662), .A1(n452), .B0(n968), .B1(n460), .Y(n1114) );
  OAI22XL U1673 ( .A0(n1662), .A1(n451), .B0(n968), .B1(n459), .Y(n1109) );
  OAI22XL U1674 ( .A0(n1662), .A1(n450), .B0(n968), .B1(n458), .Y(n1104) );
  NOR4X1 U1675 ( .A(n1688), .B(index_b[5]), .C(index_b[6]), .D(index_b[7]), 
        .Y(n1272) );
  NAND2X1 U1676 ( .A(cur_state[1]), .B(n225), .Y(n941) );
  OAI22XL U1677 ( .A0(n1815), .A1(n1594), .B0(n1634), .B1(n558), .Y(n1487) );
  CLKINVX1 U1678 ( .A(data_out_b[3]), .Y(n1815) );
  OAI22XL U1679 ( .A0(n1814), .A1(n1594), .B0(n1634), .B1(n557), .Y(n1486) );
  CLKINVX1 U1680 ( .A(data_out_b[4]), .Y(n1814) );
  OAI22XL U1681 ( .A0(n1813), .A1(n1594), .B0(n1634), .B1(n556), .Y(n1485) );
  CLKINVX1 U1682 ( .A(data_out_b[5]), .Y(n1813) );
  OAI22XL U1683 ( .A0(n1812), .A1(n1594), .B0(n1634), .B1(n555), .Y(n1484) );
  CLKINVX1 U1684 ( .A(data_out_b[6]), .Y(n1812) );
  OAI22XL U1685 ( .A0(n1811), .A1(n1594), .B0(n1634), .B1(n554), .Y(n1483) );
  CLKINVX1 U1686 ( .A(data_out_b[7]), .Y(n1811) );
  OAI22XL U1687 ( .A0(n1810), .A1(n1594), .B0(n1634), .B1(n553), .Y(n1474) );
  CLKINVX1 U1688 ( .A(data_out_b[8]), .Y(n1810) );
  OAI22XL U1689 ( .A0(n1809), .A1(n1594), .B0(n1634), .B1(n552), .Y(n1473) );
  CLKINVX1 U1690 ( .A(data_out_b[9]), .Y(n1809) );
  OAI22XL U1691 ( .A0(n1808), .A1(n1594), .B0(n1634), .B1(n551), .Y(n1472) );
  CLKINVX1 U1692 ( .A(data_out_b[10]), .Y(n1808) );
  OAI22XL U1693 ( .A0(n1807), .A1(n1594), .B0(n1634), .B1(n550), .Y(n1471) );
  CLKINVX1 U1694 ( .A(data_out_b[11]), .Y(n1807) );
  OAI22XL U1695 ( .A0(n1806), .A1(n1594), .B0(n1634), .B1(n549), .Y(n1470) );
  CLKINVX1 U1696 ( .A(data_out_b[12]), .Y(n1806) );
  OAI22XL U1697 ( .A0(n1805), .A1(n1594), .B0(n1634), .B1(n548), .Y(n1469) );
  CLKINVX1 U1698 ( .A(data_out_b[13]), .Y(n1805) );
  OAI22XL U1699 ( .A0(n1804), .A1(n1594), .B0(n1634), .B1(n547), .Y(n1468) );
  CLKINVX1 U1700 ( .A(data_out_b[14]), .Y(n1804) );
  OAI22XL U1701 ( .A0(n1803), .A1(n1594), .B0(n1634), .B1(n546), .Y(n1467) );
  CLKINVX1 U1702 ( .A(data_out_b[15]), .Y(n1803) );
  OAI22XL U1703 ( .A0(n1818), .A1(n1594), .B0(n1634), .B1(n561), .Y(n1490) );
  CLKINVX1 U1704 ( .A(data_out_b[0]), .Y(n1818) );
  OAI22XL U1705 ( .A0(n1817), .A1(n1594), .B0(n1908), .B1(n560), .Y(n1489) );
  CLKINVX1 U1706 ( .A(data_out_b[1]), .Y(n1817) );
  OAI22XL U1707 ( .A0(n1816), .A1(n1594), .B0(n1908), .B1(n559), .Y(n1488) );
  CLKINVX1 U1708 ( .A(data_out_b[2]), .Y(n1816) );
  OAI22XL U1709 ( .A0(n1850), .A1(n1645), .B0(n1648), .B1(n353), .Y(n1394) );
  CLKINVX1 U1710 ( .A(data_out_a[0]), .Y(n1850) );
  OAI22XL U1711 ( .A0(n1849), .A1(n1645), .B0(n1648), .B1(n352), .Y(n1393) );
  CLKINVX1 U1712 ( .A(data_out_a[1]), .Y(n1849) );
  OAI22XL U1713 ( .A0(n1848), .A1(n1645), .B0(n1647), .B1(n351), .Y(n1392) );
  CLKINVX1 U1714 ( .A(data_out_a[2]), .Y(n1848) );
  OAI22XL U1715 ( .A0(n1847), .A1(n1645), .B0(n1648), .B1(n350), .Y(n1391) );
  CLKINVX1 U1716 ( .A(data_out_a[3]), .Y(n1847) );
  OAI22XL U1717 ( .A0(n1846), .A1(n1645), .B0(n1647), .B1(n349), .Y(n1390) );
  CLKINVX1 U1718 ( .A(data_out_a[4]), .Y(n1846) );
  OAI22XL U1719 ( .A0(n1845), .A1(n1645), .B0(n1648), .B1(n348), .Y(n1389) );
  CLKINVX1 U1720 ( .A(data_out_a[5]), .Y(n1845) );
  OAI22XL U1721 ( .A0(n1844), .A1(n1645), .B0(n1647), .B1(n347), .Y(n1388) );
  CLKINVX1 U1722 ( .A(data_out_a[6]), .Y(n1844) );
  OAI22XL U1723 ( .A0(n1843), .A1(n1645), .B0(n1510), .B1(n346), .Y(n1387) );
  CLKINVX1 U1724 ( .A(data_out_a[7]), .Y(n1843) );
  OAI22XL U1725 ( .A0(n1842), .A1(n1645), .B0(n1510), .B1(n345), .Y(n1386) );
  CLKINVX1 U1726 ( .A(n1578), .Y(n1842) );
  OAI22XL U1727 ( .A0(n1841), .A1(n1645), .B0(n1648), .B1(n344), .Y(n1385) );
  CLKINVX1 U1728 ( .A(n1579), .Y(n1841) );
  OAI22XL U1729 ( .A0(n1840), .A1(n1645), .B0(n1647), .B1(n343), .Y(n1384) );
  CLKINVX1 U1730 ( .A(n1580), .Y(n1840) );
  OAI22XL U1731 ( .A0(n1839), .A1(n1645), .B0(n1647), .B1(n342), .Y(n1383) );
  CLKINVX1 U1732 ( .A(n1581), .Y(n1839) );
  OAI22XL U1733 ( .A0(n1838), .A1(n1646), .B0(n1647), .B1(n341), .Y(n1382) );
  CLKINVX1 U1734 ( .A(n1582), .Y(n1838) );
  OAI22XL U1735 ( .A0(n1837), .A1(n1646), .B0(n1647), .B1(n340), .Y(n1381) );
  CLKINVX1 U1736 ( .A(n1583), .Y(n1837) );
  OAI22XL U1737 ( .A0(n1836), .A1(n1646), .B0(n1647), .B1(n339), .Y(n1380) );
  CLKINVX1 U1738 ( .A(n1584), .Y(n1836) );
  OAI22XL U1739 ( .A0(n1835), .A1(n1646), .B0(n1647), .B1(n338), .Y(n1379) );
  CLKINVX1 U1740 ( .A(n1585), .Y(n1835) );
  OAI22XL U1741 ( .A0(n1834), .A1(n1646), .B0(n1647), .B1(n337), .Y(n1378) );
  CLKINVX1 U1742 ( .A(n1586), .Y(n1834) );
  OAI22XL U1743 ( .A0(n1833), .A1(n1646), .B0(n1647), .B1(n336), .Y(n1377) );
  CLKINVX1 U1744 ( .A(n1587), .Y(n1833) );
  OAI22XL U1745 ( .A0(n1832), .A1(n1646), .B0(n1647), .B1(n335), .Y(n1376) );
  CLKINVX1 U1746 ( .A(n1588), .Y(n1832) );
  OAI22XL U1747 ( .A0(n1831), .A1(n1646), .B0(n1648), .B1(n334), .Y(n1375) );
  CLKINVX1 U1748 ( .A(n1589), .Y(n1831) );
  OAI22XL U1749 ( .A0(n1830), .A1(n1646), .B0(n1647), .B1(n333), .Y(n1374) );
  CLKINVX1 U1750 ( .A(n1590), .Y(n1830) );
  OAI22XL U1751 ( .A0(n1829), .A1(n1646), .B0(n1648), .B1(n332), .Y(n1373) );
  CLKINVX1 U1752 ( .A(n1591), .Y(n1829) );
  OAI22XL U1753 ( .A0(n1828), .A1(n1646), .B0(n1647), .B1(n331), .Y(n1372) );
  CLKINVX1 U1754 ( .A(n1592), .Y(n1828) );
  OAI22XL U1755 ( .A0(n1827), .A1(n1646), .B0(n1648), .B1(n330), .Y(n1371) );
  CLKINVX1 U1756 ( .A(n1593), .Y(n1827) );
  OAI22XL U1757 ( .A0(n1826), .A1(n1645), .B0(n1647), .B1(n329), .Y(n1370) );
  CLKINVX1 U1758 ( .A(data_out_a[24]), .Y(n1826) );
  OAI22XL U1759 ( .A0(n1825), .A1(n1646), .B0(n1648), .B1(n328), .Y(n1369) );
  CLKINVX1 U1760 ( .A(data_out_a[25]), .Y(n1825) );
  OAI22XL U1761 ( .A0(n1824), .A1(n1645), .B0(n1648), .B1(n327), .Y(n1368) );
  CLKINVX1 U1762 ( .A(data_out_a[26]), .Y(n1824) );
  OAI22XL U1763 ( .A0(n1823), .A1(n1646), .B0(n1648), .B1(n326), .Y(n1367) );
  CLKINVX1 U1764 ( .A(data_out_a[27]), .Y(n1823) );
  OAI22XL U1765 ( .A0(n1822), .A1(n1645), .B0(n1648), .B1(n325), .Y(n1366) );
  CLKINVX1 U1766 ( .A(data_out_a[28]), .Y(n1822) );
  OAI22XL U1767 ( .A0(n1821), .A1(n1646), .B0(n1648), .B1(n324), .Y(n1365) );
  CLKINVX1 U1768 ( .A(data_out_a[29]), .Y(n1821) );
  OAI22XL U1769 ( .A0(n1820), .A1(n1645), .B0(n1648), .B1(n323), .Y(n1364) );
  CLKINVX1 U1770 ( .A(data_out_a[30]), .Y(n1820) );
  OAI22XL U1771 ( .A0(n1819), .A1(n1646), .B0(n1648), .B1(n322), .Y(n1363) );
  CLKINVX1 U1772 ( .A(data_out_a[31]), .Y(n1819) );
  OAI211X1 U1773 ( .A0(n1786), .A1(n1675), .B0(n901), .C0(n902), .Y(n900) );
  NAND2X1 U1774 ( .A(w23[0]), .B(n1672), .Y(n901) );
  AOI22X1 U1775 ( .A0(w22[0]), .A1(n1678), .B0(w21[0]), .B1(n1676), .Y(n902)
         );
  OAI211X1 U1776 ( .A0(n1770), .A1(n1675), .B0(n955), .C0(n956), .Y(n954) );
  NAND2X1 U1777 ( .A(w13[0]), .B(n1672), .Y(n955) );
  AOI22X1 U1778 ( .A0(w12[0]), .A1(n1678), .B0(w11[0]), .B1(n1676), .Y(n956)
         );
  CLKBUFX3 U1779 ( .A(n969), .Y(n1655) );
  NAND3X1 U1780 ( .A(n1629), .B(n700), .C(n1225), .Y(n969) );
  OAI2BB2XL U1781 ( .B0(n1608), .B1(n1175), .A0N(b21[0]), .A1N(n1608), .Y(
        n1410) );
  AOI222XL U1782 ( .A0(\matrix_b[5][24] ), .A1(n1668), .B0(\matrix_b[0][16] ), 
        .B1(n1909), .C0(\matrix_b[8][16] ), .C1(n1651), .Y(n1175) );
  OAI2BB2XL U1783 ( .B0(n1608), .B1(n1172), .A0N(b21[3]), .A1N(n1608), .Y(
        n1407) );
  AOI222XL U1784 ( .A0(\matrix_b[5][27] ), .A1(n1668), .B0(\matrix_b[0][19] ), 
        .B1(n1909), .C0(\matrix_b[8][19] ), .C1(n1651), .Y(n1172) );
  OAI2BB2XL U1785 ( .B0(n1608), .B1(n1171), .A0N(b21[4]), .A1N(n1608), .Y(
        n1406) );
  AOI222XL U1786 ( .A0(\matrix_b[5][28] ), .A1(n1668), .B0(\matrix_b[0][20] ), 
        .B1(n1909), .C0(\matrix_b[8][20] ), .C1(n1651), .Y(n1171) );
  OAI2BB2XL U1787 ( .B0(n1608), .B1(n1170), .A0N(b21[5]), .A1N(n1608), .Y(
        n1405) );
  AOI222XL U1788 ( .A0(\matrix_b[5][29] ), .A1(n1668), .B0(\matrix_b[0][21] ), 
        .B1(n1909), .C0(\matrix_b[8][21] ), .C1(n1651), .Y(n1170) );
  OAI2BB2XL U1789 ( .B0(n1608), .B1(n1169), .A0N(b21[6]), .A1N(n1608), .Y(
        n1404) );
  AOI222XL U1790 ( .A0(\matrix_b[5][30] ), .A1(n1668), .B0(\matrix_b[0][22] ), 
        .B1(n1909), .C0(\matrix_b[8][22] ), .C1(n1651), .Y(n1169) );
  OAI2BB2XL U1791 ( .B0(n1608), .B1(n1168), .A0N(b21[7]), .A1N(n1608), .Y(
        n1403) );
  AOI222XL U1792 ( .A0(\matrix_b[5][31] ), .A1(n1668), .B0(\matrix_b[0][23] ), 
        .B1(n1909), .C0(\matrix_b[8][23] ), .C1(n1651), .Y(n1168) );
  OAI2BB2XL U1793 ( .B0(n1609), .B1(n1162), .A0N(b11[0]), .A1N(n1609), .Y(
        n1402) );
  AOI222XL U1794 ( .A0(\matrix_b[4][24] ), .A1(n1671), .B0(\matrix_b[0][24] ), 
        .B1(n1912), .C0(\matrix_b[8][24] ), .C1(n1660), .Y(n1162) );
  OAI2BB2XL U1795 ( .B0(n1609), .B1(n1161), .A0N(b11[1]), .A1N(n1609), .Y(
        n1401) );
  AOI222XL U1796 ( .A0(\matrix_b[4][25] ), .A1(n1671), .B0(\matrix_b[0][25] ), 
        .B1(n1912), .C0(\matrix_b[8][25] ), .C1(n1660), .Y(n1161) );
  OAI2BB2XL U1797 ( .B0(n1609), .B1(n1160), .A0N(b11[2]), .A1N(n1609), .Y(
        n1400) );
  AOI222XL U1798 ( .A0(\matrix_b[4][26] ), .A1(n1671), .B0(\matrix_b[0][26] ), 
        .B1(n1912), .C0(\matrix_b[8][26] ), .C1(n1660), .Y(n1160) );
  OAI2BB2XL U1799 ( .B0(n1609), .B1(n1159), .A0N(b11[3]), .A1N(n1609), .Y(
        n1399) );
  AOI222XL U1800 ( .A0(\matrix_b[4][27] ), .A1(n1671), .B0(\matrix_b[0][27] ), 
        .B1(n1912), .C0(\matrix_b[8][27] ), .C1(n1660), .Y(n1159) );
  OAI2BB2XL U1801 ( .B0(n1609), .B1(n1158), .A0N(b11[4]), .A1N(n1609), .Y(
        n1398) );
  AOI222XL U1802 ( .A0(\matrix_b[4][28] ), .A1(n1671), .B0(\matrix_b[0][28] ), 
        .B1(n1912), .C0(\matrix_b[8][28] ), .C1(n1660), .Y(n1158) );
  OAI2BB2XL U1803 ( .B0(n1609), .B1(n1157), .A0N(b11[5]), .A1N(n1609), .Y(
        n1397) );
  AOI222XL U1804 ( .A0(\matrix_b[4][29] ), .A1(n1671), .B0(\matrix_b[0][29] ), 
        .B1(n1912), .C0(\matrix_b[8][29] ), .C1(n1660), .Y(n1157) );
  OAI2BB2XL U1805 ( .B0(n1609), .B1(n1156), .A0N(b11[6]), .A1N(n1609), .Y(
        n1396) );
  AOI222XL U1806 ( .A0(\matrix_b[4][30] ), .A1(n1671), .B0(\matrix_b[0][30] ), 
        .B1(n1912), .C0(\matrix_b[8][30] ), .C1(n1660), .Y(n1156) );
  OAI2BB2XL U1807 ( .B0(n1609), .B1(n1155), .A0N(b11[7]), .A1N(n1609), .Y(
        n1395) );
  AOI222XL U1808 ( .A0(\matrix_b[4][31] ), .A1(n1671), .B0(\matrix_b[0][31] ), 
        .B1(n1912), .C0(\matrix_b[8][31] ), .C1(n1660), .Y(n1155) );
  OAI2BB2XL U1809 ( .B0(n1606), .B1(n1195), .A0N(b41[0]), .A1N(n1606), .Y(
        n1426) );
  AOI222XL U1810 ( .A0(\matrix_b[0][0] ), .A1(n1571), .B0(n1910), .B1(
        \matrix_b[8][0] ), .C0(\matrix_b[7][24] ), .C1(n1663), .Y(n1195) );
  OAI2BB2XL U1811 ( .B0(n1606), .B1(n1194), .A0N(b41[1]), .A1N(n1606), .Y(
        n1425) );
  AOI222XL U1812 ( .A0(\matrix_b[0][1] ), .A1(n1571), .B0(n1910), .B1(
        \matrix_b[8][1] ), .C0(\matrix_b[7][25] ), .C1(n1663), .Y(n1194) );
  OAI2BB2XL U1813 ( .B0(n1606), .B1(n1193), .A0N(b41[2]), .A1N(n1606), .Y(
        n1424) );
  AOI222XL U1814 ( .A0(\matrix_b[0][2] ), .A1(n1571), .B0(n1910), .B1(
        \matrix_b[8][2] ), .C0(\matrix_b[7][26] ), .C1(n1663), .Y(n1193) );
  OAI2BB2XL U1815 ( .B0(n1606), .B1(n1192), .A0N(b41[3]), .A1N(n1606), .Y(
        n1423) );
  AOI222XL U1816 ( .A0(\matrix_b[0][3] ), .A1(n1571), .B0(n1910), .B1(
        \matrix_b[8][3] ), .C0(\matrix_b[7][27] ), .C1(n1663), .Y(n1192) );
  OAI2BB2XL U1817 ( .B0(n1606), .B1(n1191), .A0N(b41[4]), .A1N(n1606), .Y(
        n1422) );
  AOI222XL U1818 ( .A0(\matrix_b[0][4] ), .A1(n1571), .B0(n1910), .B1(
        \matrix_b[8][4] ), .C0(\matrix_b[7][28] ), .C1(n1663), .Y(n1191) );
  OAI2BB2XL U1819 ( .B0(n1606), .B1(n1190), .A0N(b41[5]), .A1N(n1606), .Y(
        n1421) );
  AOI222XL U1820 ( .A0(\matrix_b[0][5] ), .A1(n1571), .B0(n1910), .B1(
        \matrix_b[8][5] ), .C0(\matrix_b[7][29] ), .C1(n1663), .Y(n1190) );
  OAI2BB2XL U1821 ( .B0(n1606), .B1(n1189), .A0N(b41[6]), .A1N(n1606), .Y(
        n1420) );
  AOI222XL U1822 ( .A0(\matrix_b[0][6] ), .A1(n1571), .B0(n1910), .B1(
        \matrix_b[8][6] ), .C0(\matrix_b[7][30] ), .C1(n1663), .Y(n1189) );
  OAI2BB2XL U1823 ( .B0(n1606), .B1(n1188), .A0N(b41[7]), .A1N(n1606), .Y(
        n1419) );
  AOI222XL U1824 ( .A0(\matrix_b[0][7] ), .A1(n1571), .B0(n1910), .B1(
        \matrix_b[8][7] ), .C0(\matrix_b[7][31] ), .C1(n1663), .Y(n1188) );
  OAI2BB2XL U1825 ( .B0(n1607), .B1(n1185), .A0N(b31[0]), .A1N(n1607), .Y(
        n1418) );
  AOI222XL U1826 ( .A0(\matrix_b[6][24] ), .A1(n1657), .B0(\matrix_b[0][8] ), 
        .B1(n1654), .C0(n1911), .C1(\matrix_b[8][8] ), .Y(n1185) );
  OAI2BB2XL U1827 ( .B0(n1607), .B1(n1184), .A0N(b31[1]), .A1N(n1607), .Y(
        n1417) );
  AOI222XL U1828 ( .A0(\matrix_b[6][25] ), .A1(n1657), .B0(\matrix_b[0][9] ), 
        .B1(n1654), .C0(n1911), .C1(\matrix_b[8][9] ), .Y(n1184) );
  OAI2BB2XL U1829 ( .B0(n1607), .B1(n1183), .A0N(b31[2]), .A1N(n1607), .Y(
        n1416) );
  AOI222XL U1830 ( .A0(\matrix_b[6][26] ), .A1(n1657), .B0(\matrix_b[0][10] ), 
        .B1(n1654), .C0(n1911), .C1(\matrix_b[8][10] ), .Y(n1183) );
  OAI2BB2XL U1831 ( .B0(n1607), .B1(n1182), .A0N(b31[3]), .A1N(n1607), .Y(
        n1415) );
  AOI222XL U1832 ( .A0(\matrix_b[6][27] ), .A1(n1657), .B0(\matrix_b[0][11] ), 
        .B1(n1654), .C0(n1911), .C1(\matrix_b[8][11] ), .Y(n1182) );
  OAI2BB2XL U1833 ( .B0(n1607), .B1(n1181), .A0N(b31[4]), .A1N(n1607), .Y(
        n1414) );
  AOI222XL U1834 ( .A0(\matrix_b[6][28] ), .A1(n1657), .B0(\matrix_b[0][12] ), 
        .B1(n1653), .C0(n1911), .C1(\matrix_b[8][12] ), .Y(n1181) );
  OAI2BB2XL U1835 ( .B0(n1607), .B1(n1180), .A0N(b31[5]), .A1N(n1607), .Y(
        n1413) );
  AOI222XL U1836 ( .A0(\matrix_b[6][29] ), .A1(n1657), .B0(\matrix_b[0][13] ), 
        .B1(n1653), .C0(\matrix_b[8][13] ), .C1(n1911), .Y(n1180) );
  OAI2BB2XL U1837 ( .B0(n1607), .B1(n1179), .A0N(b31[6]), .A1N(n1607), .Y(
        n1412) );
  AOI222XL U1838 ( .A0(\matrix_b[6][30] ), .A1(n1657), .B0(\matrix_b[0][14] ), 
        .B1(n1654), .C0(\matrix_b[8][14] ), .C1(n1911), .Y(n1179) );
  OAI2BB2XL U1839 ( .B0(n1607), .B1(n1178), .A0N(b31[7]), .A1N(n1607), .Y(
        n1411) );
  AOI222XL U1840 ( .A0(\matrix_b[6][31] ), .A1(n1657), .B0(\matrix_b[0][15] ), 
        .B1(n1653), .C0(\matrix_b[8][15] ), .C1(n1911), .Y(n1178) );
  OAI2BB2XL U1841 ( .B0(n1608), .B1(n1174), .A0N(b21[1]), .A1N(n1608), .Y(
        n1409) );
  AOI222XL U1842 ( .A0(\matrix_b[5][25] ), .A1(n1668), .B0(\matrix_b[0][17] ), 
        .B1(n1909), .C0(\matrix_b[8][17] ), .C1(n1650), .Y(n1174) );
  OAI2BB2XL U1843 ( .B0(n1608), .B1(n1173), .A0N(b21[2]), .A1N(n1608), .Y(
        n1408) );
  AOI222XL U1844 ( .A0(\matrix_b[5][26] ), .A1(n1668), .B0(\matrix_b[0][18] ), 
        .B1(n1909), .C0(\matrix_b[8][18] ), .C1(n1650), .Y(n1173) );
  OAI2BB2XL U1845 ( .B0(n1006), .B1(n1613), .A0N(a11[0]), .A1N(n1613), .Y(
        n1338) );
  NOR4X1 U1846 ( .A(n1009), .B(n1010), .C(n1011), .D(n1012), .Y(n1006) );
  OAI222XL U1847 ( .A0(n973), .A1(n233), .B0(n974), .B1(n513), .C0(n1604), 
        .C1(n241), .Y(n1009) );
  OAI222XL U1848 ( .A0(n1595), .A1(n505), .B0(n1652), .B1(n249), .C0(n1649), 
        .C1(n497), .Y(n1010) );
  OAI2BB2XL U1849 ( .B0(n1001), .B1(n1613), .A0N(a11[1]), .A1N(n1613), .Y(
        n1337) );
  NOR4X1 U1850 ( .A(n1002), .B(n1003), .C(n1004), .D(n1005), .Y(n1001) );
  OAI222XL U1851 ( .A0(n973), .A1(n232), .B0(n974), .B1(n512), .C0(n1604), 
        .C1(n240), .Y(n1002) );
  OAI222XL U1852 ( .A0(n1595), .A1(n504), .B0(n1652), .B1(n248), .C0(n1649), 
        .C1(n496), .Y(n1003) );
  OAI2BB2XL U1853 ( .B0(n996), .B1(n1613), .A0N(a11[2]), .A1N(n1613), .Y(n1336) );
  NOR4X1 U1854 ( .A(n997), .B(n998), .C(n999), .D(n1000), .Y(n996) );
  OAI222XL U1855 ( .A0(n973), .A1(n231), .B0(n974), .B1(n511), .C0(n1604), 
        .C1(n239), .Y(n997) );
  OAI222XL U1856 ( .A0(n1595), .A1(n503), .B0(n1652), .B1(n247), .C0(n972), 
        .C1(n495), .Y(n998) );
  OAI2BB2XL U1857 ( .B0(n991), .B1(n1613), .A0N(a11[3]), .A1N(n1613), .Y(n1335) );
  NOR4X1 U1858 ( .A(n992), .B(n993), .C(n994), .D(n995), .Y(n991) );
  OAI222XL U1859 ( .A0(n973), .A1(n230), .B0(n974), .B1(n510), .C0(n1604), 
        .C1(n238), .Y(n992) );
  OAI222XL U1860 ( .A0(n1595), .A1(n502), .B0(n1652), .B1(n246), .C0(n972), 
        .C1(n494), .Y(n993) );
  OAI2BB2XL U1861 ( .B0(n986), .B1(n1613), .A0N(a11[4]), .A1N(n1613), .Y(n1334) );
  NOR4X1 U1862 ( .A(n987), .B(n988), .C(n989), .D(n990), .Y(n986) );
  OAI222XL U1863 ( .A0(n973), .A1(n229), .B0(n974), .B1(n509), .C0(n1604), 
        .C1(n237), .Y(n987) );
  OAI222XL U1864 ( .A0(n1662), .A1(n381), .B0(n1659), .B1(n485), .C0(n1656), 
        .C1(n373), .Y(n989) );
  OAI2BB2XL U1865 ( .B0(n981), .B1(n1613), .A0N(a11[5]), .A1N(n1613), .Y(n1333) );
  NOR4X1 U1866 ( .A(n982), .B(n983), .C(n984), .D(n985), .Y(n981) );
  OAI222XL U1867 ( .A0(n973), .A1(n228), .B0(n974), .B1(n508), .C0(n1604), 
        .C1(n236), .Y(n982) );
  OAI222XL U1868 ( .A0(n1662), .A1(n380), .B0(n1659), .B1(n484), .C0(n1655), 
        .C1(n372), .Y(n984) );
  OAI2BB2XL U1869 ( .B0(n976), .B1(n1613), .A0N(a11[6]), .A1N(n1613), .Y(n1332) );
  NOR4X1 U1870 ( .A(n977), .B(n978), .C(n979), .D(n980), .Y(n976) );
  OAI222XL U1871 ( .A0(n973), .A1(n227), .B0(n974), .B1(n507), .C0(n1604), 
        .C1(n235), .Y(n977) );
  OAI222XL U1872 ( .A0(n1662), .A1(n379), .B0(n1659), .B1(n483), .C0(n1655), 
        .C1(n371), .Y(n979) );
  OAI2BB2XL U1873 ( .B0(n958), .B1(n1613), .A0N(a11[7]), .A1N(n1613), .Y(n1331) );
  NOR4X1 U1874 ( .A(n960), .B(n961), .C(n962), .D(n963), .Y(n958) );
  OAI222XL U1875 ( .A0(n973), .A1(n226), .B0(n974), .B1(n506), .C0(n1604), 
        .C1(n234), .Y(n960) );
  OAI222XL U1876 ( .A0(n1662), .A1(n378), .B0(n1659), .B1(n482), .C0(n1655), 
        .C1(n370), .Y(n962) );
  OAI2BB2XL U1877 ( .B0(n1095), .B1(n1611), .A0N(a13[0]), .A1N(n1611), .Y(
        n1354) );
  NOR4X1 U1878 ( .A(n1096), .B(n1097), .C(n1098), .D(n1099), .Y(n1095) );
  OAI22XL U1879 ( .A0(n1649), .A1(n449), .B0(n1652), .B1(n297), .Y(n1096) );
  OAI22XL U1880 ( .A0(n1666), .A1(n321), .B0(n1656), .B1(n425), .Y(n1098) );
  OAI2BB2XL U1881 ( .B0(n1090), .B1(n1611), .A0N(a13[1]), .A1N(n1611), .Y(
        n1353) );
  NOR4X1 U1882 ( .A(n1091), .B(n1092), .C(n1093), .D(n1094), .Y(n1090) );
  OAI22XL U1883 ( .A0(n1649), .A1(n448), .B0(n1652), .B1(n296), .Y(n1091) );
  OAI22XL U1884 ( .A0(n1666), .A1(n320), .B0(n1655), .B1(n424), .Y(n1093) );
  OAI2BB2XL U1885 ( .B0(n1085), .B1(n1611), .A0N(a13[2]), .A1N(n1611), .Y(
        n1352) );
  NOR4X1 U1886 ( .A(n1086), .B(n1087), .C(n1088), .D(n1089), .Y(n1085) );
  OAI22XL U1887 ( .A0(n1649), .A1(n447), .B0(n1652), .B1(n295), .Y(n1086) );
  OAI22XL U1888 ( .A0(n1666), .A1(n319), .B0(n1655), .B1(n423), .Y(n1088) );
  OAI2BB2XL U1889 ( .B0(n1080), .B1(n1611), .A0N(a13[3]), .A1N(n1611), .Y(
        n1351) );
  NOR4X1 U1890 ( .A(n1081), .B(n1082), .C(n1083), .D(n1084), .Y(n1080) );
  OAI22XL U1891 ( .A0(n1649), .A1(n446), .B0(n1652), .B1(n294), .Y(n1081) );
  OAI22XL U1892 ( .A0(n1666), .A1(n318), .B0(n1655), .B1(n422), .Y(n1083) );
  OAI2BB2XL U1893 ( .B0(n1075), .B1(n1611), .A0N(a13[4]), .A1N(n1611), .Y(
        n1350) );
  NOR4X1 U1894 ( .A(n1076), .B(n1077), .C(n1078), .D(n1079), .Y(n1075) );
  OAI22XL U1895 ( .A0(n1649), .A1(n445), .B0(n1652), .B1(n293), .Y(n1076) );
  OAI22XL U1896 ( .A0(n1666), .A1(n317), .B0(n1656), .B1(n421), .Y(n1078) );
  OAI2BB2XL U1897 ( .B0(n1070), .B1(n1611), .A0N(a13[5]), .A1N(n1611), .Y(
        n1349) );
  NOR4X1 U1898 ( .A(n1071), .B(n1072), .C(n1073), .D(n1074), .Y(n1070) );
  OAI22XL U1899 ( .A0(n1649), .A1(n444), .B0(n1652), .B1(n292), .Y(n1071) );
  OAI22XL U1900 ( .A0(n1667), .A1(n316), .B0(n1656), .B1(n420), .Y(n1073) );
  OAI2BB2XL U1901 ( .B0(n1065), .B1(n1611), .A0N(a13[6]), .A1N(n1611), .Y(
        n1348) );
  NOR4X1 U1902 ( .A(n1066), .B(n1067), .C(n1068), .D(n1069), .Y(n1065) );
  OAI22XL U1903 ( .A0(n1649), .A1(n443), .B0(n1652), .B1(n291), .Y(n1066) );
  OAI22XL U1904 ( .A0(n965), .A1(n315), .B0(n1656), .B1(n419), .Y(n1068) );
  OAI2BB2XL U1905 ( .B0(n1059), .B1(n1611), .A0N(a13[7]), .A1N(n1611), .Y(
        n1347) );
  NOR4X1 U1906 ( .A(n1061), .B(n1062), .C(n1063), .D(n1064), .Y(n1059) );
  OAI22XL U1907 ( .A0(n1649), .A1(n442), .B0(n1652), .B1(n290), .Y(n1061) );
  OAI22XL U1908 ( .A0(n965), .A1(n314), .B0(n1656), .B1(n418), .Y(n1063) );
  OAI2BB2XL U1909 ( .B0(n1137), .B1(n1610), .A0N(a14[0]), .A1N(n1610), .Y(
        n1362) );
  NOR4X1 U1910 ( .A(n1141), .B(n1142), .C(n1143), .D(n1144), .Y(n1137) );
  OAI22XL U1911 ( .A0(n972), .A1(n473), .B0(n1595), .B1(n481), .Y(n1141) );
  OAI22XL U1912 ( .A0(n1666), .A1(n345), .B0(n1655), .B1(n353), .Y(n1143) );
  OAI2BB2XL U1913 ( .B0(n1132), .B1(n1610), .A0N(a14[1]), .A1N(n1610), .Y(
        n1361) );
  NOR4X1 U1914 ( .A(n1133), .B(n1134), .C(n1135), .D(n1136), .Y(n1132) );
  OAI22XL U1915 ( .A0(n972), .A1(n472), .B0(n1595), .B1(n480), .Y(n1133) );
  OAI22XL U1916 ( .A0(n1666), .A1(n344), .B0(n1655), .B1(n352), .Y(n1135) );
  OAI2BB2XL U1917 ( .B0(n1127), .B1(n1610), .A0N(a14[2]), .A1N(n1610), .Y(
        n1360) );
  NOR4X1 U1918 ( .A(n1128), .B(n1129), .C(n1130), .D(n1131), .Y(n1127) );
  OAI22XL U1919 ( .A0(n972), .A1(n471), .B0(n1595), .B1(n479), .Y(n1128) );
  OAI22XL U1920 ( .A0(n1666), .A1(n343), .B0(n1655), .B1(n351), .Y(n1130) );
  OAI2BB2XL U1921 ( .B0(n1122), .B1(n1610), .A0N(a14[3]), .A1N(n1610), .Y(
        n1359) );
  NOR4X1 U1922 ( .A(n1123), .B(n1124), .C(n1125), .D(n1126), .Y(n1122) );
  OAI22XL U1923 ( .A0(n1649), .A1(n470), .B0(n1595), .B1(n478), .Y(n1123) );
  OAI22XL U1924 ( .A0(n1666), .A1(n342), .B0(n1655), .B1(n350), .Y(n1125) );
  OAI2BB2XL U1925 ( .B0(n1117), .B1(n1610), .A0N(a14[4]), .A1N(n1610), .Y(
        n1358) );
  NOR4X1 U1926 ( .A(n1118), .B(n1119), .C(n1120), .D(n1121), .Y(n1117) );
  OAI22XL U1927 ( .A0(n1649), .A1(n469), .B0(n1595), .B1(n477), .Y(n1118) );
  OAI22XL U1928 ( .A0(n1666), .A1(n341), .B0(n1655), .B1(n349), .Y(n1120) );
  OAI2BB2XL U1929 ( .B0(n1112), .B1(n1610), .A0N(a14[5]), .A1N(n1610), .Y(
        n1357) );
  NOR4X1 U1930 ( .A(n1113), .B(n1114), .C(n1115), .D(n1116), .Y(n1112) );
  OAI22XL U1931 ( .A0(n1649), .A1(n468), .B0(n1595), .B1(n476), .Y(n1113) );
  OAI22XL U1932 ( .A0(n1666), .A1(n340), .B0(n969), .B1(n348), .Y(n1115) );
  OAI2BB2XL U1933 ( .B0(n1107), .B1(n1610), .A0N(a14[6]), .A1N(n1610), .Y(
        n1356) );
  NOR4X1 U1934 ( .A(n1108), .B(n1109), .C(n1110), .D(n1111), .Y(n1107) );
  OAI22XL U1935 ( .A0(n1649), .A1(n467), .B0(n1595), .B1(n475), .Y(n1108) );
  OAI22XL U1936 ( .A0(n1666), .A1(n339), .B0(n969), .B1(n347), .Y(n1110) );
  OAI2BB2XL U1937 ( .B0(n1101), .B1(n1610), .A0N(a14[7]), .A1N(n1610), .Y(
        n1355) );
  NOR4X1 U1938 ( .A(n1103), .B(n1104), .C(n1105), .D(n1106), .Y(n1101) );
  OAI22XL U1939 ( .A0(n1649), .A1(n466), .B0(n1595), .B1(n474), .Y(n1103) );
  OAI22XL U1940 ( .A0(n1666), .A1(n338), .B0(n969), .B1(n346), .Y(n1105) );
  OAI2BB2XL U1941 ( .B0(n1051), .B1(n1612), .A0N(a12[0]), .A1N(n1612), .Y(
        n1346) );
  NOR4X1 U1942 ( .A(n1053), .B(n1054), .C(n1055), .D(n1056), .Y(n1051) );
  OAI22XL U1943 ( .A0(n1652), .A1(n273), .B0(n1604), .B1(n265), .Y(n1053) );
  OAI22XL U1944 ( .A0(n965), .A1(n393), .B0(n1656), .B1(n401), .Y(n1055) );
  OAI2BB2XL U1945 ( .B0(n1046), .B1(n1612), .A0N(a12[1]), .A1N(n1612), .Y(
        n1345) );
  NOR4X1 U1946 ( .A(n1047), .B(n1048), .C(n1049), .D(n1050), .Y(n1046) );
  OAI22XL U1947 ( .A0(n1652), .A1(n272), .B0(n1604), .B1(n264), .Y(n1047) );
  OAI22XL U1948 ( .A0(n1666), .A1(n392), .B0(n1656), .B1(n400), .Y(n1049) );
  OAI2BB2XL U1949 ( .B0(n1041), .B1(n1612), .A0N(a12[2]), .A1N(n1612), .Y(
        n1344) );
  NOR4X1 U1950 ( .A(n1042), .B(n1043), .C(n1044), .D(n1045), .Y(n1041) );
  OAI22XL U1951 ( .A0(n1652), .A1(n271), .B0(n1604), .B1(n263), .Y(n1042) );
  OAI22XL U1952 ( .A0(n1666), .A1(n391), .B0(n1656), .B1(n399), .Y(n1044) );
  OAI2BB2XL U1953 ( .B0(n1036), .B1(n1612), .A0N(a12[3]), .A1N(n1612), .Y(
        n1343) );
  NOR4X1 U1954 ( .A(n1037), .B(n1038), .C(n1039), .D(n1040), .Y(n1036) );
  OAI22XL U1955 ( .A0(n1652), .A1(n270), .B0(n1604), .B1(n262), .Y(n1037) );
  OAI22XL U1956 ( .A0(n1666), .A1(n390), .B0(n1656), .B1(n398), .Y(n1039) );
  OAI2BB2XL U1957 ( .B0(n1031), .B1(n1612), .A0N(a12[4]), .A1N(n1612), .Y(
        n1342) );
  NOR4X1 U1958 ( .A(n1032), .B(n1033), .C(n1034), .D(n1035), .Y(n1031) );
  OAI22XL U1959 ( .A0(n971), .A1(n269), .B0(n1604), .B1(n261), .Y(n1032) );
  OAI22XL U1960 ( .A0(n1666), .A1(n389), .B0(n1656), .B1(n397), .Y(n1034) );
  OAI2BB2XL U1961 ( .B0(n1026), .B1(n1612), .A0N(a12[5]), .A1N(n1612), .Y(
        n1341) );
  NOR4X1 U1962 ( .A(n1027), .B(n1028), .C(n1029), .D(n1030), .Y(n1026) );
  OAI22XL U1963 ( .A0(n971), .A1(n268), .B0(n1604), .B1(n260), .Y(n1027) );
  OAI22XL U1964 ( .A0(n1666), .A1(n388), .B0(n1656), .B1(n396), .Y(n1029) );
  OAI2BB2XL U1965 ( .B0(n1021), .B1(n1612), .A0N(a12[6]), .A1N(n1612), .Y(
        n1340) );
  NOR4X1 U1966 ( .A(n1022), .B(n1023), .C(n1024), .D(n1025), .Y(n1021) );
  OAI22XL U1967 ( .A0(n971), .A1(n267), .B0(n1604), .B1(n259), .Y(n1022) );
  OAI22XL U1968 ( .A0(n1666), .A1(n387), .B0(n1656), .B1(n395), .Y(n1024) );
  OAI2BB2XL U1969 ( .B0(n1015), .B1(n1612), .A0N(a12[7]), .A1N(n1612), .Y(
        n1339) );
  NOR4X1 U1970 ( .A(n1017), .B(n1018), .C(n1019), .D(n1020), .Y(n1015) );
  OAI22XL U1971 ( .A0(n971), .A1(n266), .B0(n1604), .B1(n258), .Y(n1017) );
  OAI22XL U1972 ( .A0(n965), .A1(n386), .B0(n1656), .B1(n394), .Y(n1019) );
  CLKINVX1 U1973 ( .A(w44[0]), .Y(n1802) );
  CLKINVX1 U1974 ( .A(w44[1]), .Y(n1801) );
  CLKINVX1 U1975 ( .A(w44[2]), .Y(n1800) );
  CLKINVX1 U1976 ( .A(w44[3]), .Y(n1799) );
  CLKINVX1 U1977 ( .A(n1242), .Y(n1866) );
  AOI222XL U1978 ( .A0(b33[0]), .A1(n1643), .B0(\matrix_b[6][8] ), .B1(n1638), 
        .C0(\matrix_b[2][8] ), .C1(n1637), .Y(n1242) );
  CLKINVX1 U1979 ( .A(n1241), .Y(n1867) );
  AOI222XL U1980 ( .A0(b33[1]), .A1(n1643), .B0(\matrix_b[6][9] ), .B1(n1638), 
        .C0(\matrix_b[2][9] ), .C1(n1637), .Y(n1241) );
  CLKINVX1 U1981 ( .A(n1240), .Y(n1868) );
  AOI222XL U1982 ( .A0(b33[2]), .A1(n1643), .B0(\matrix_b[6][10] ), .B1(n1638), 
        .C0(\matrix_b[2][10] ), .C1(n1637), .Y(n1240) );
  CLKINVX1 U1983 ( .A(n1239), .Y(n1869) );
  AOI222XL U1984 ( .A0(b33[3]), .A1(n1643), .B0(\matrix_b[6][11] ), .B1(n1638), 
        .C0(\matrix_b[2][11] ), .C1(n1637), .Y(n1239) );
  CLKINVX1 U1985 ( .A(n1238), .Y(n1870) );
  AOI222XL U1986 ( .A0(b33[4]), .A1(n1643), .B0(\matrix_b[6][12] ), .B1(n1638), 
        .C0(\matrix_b[2][12] ), .C1(n1637), .Y(n1238) );
  CLKINVX1 U1987 ( .A(n1237), .Y(n1871) );
  AOI222XL U1988 ( .A0(b33[5]), .A1(n1643), .B0(\matrix_b[6][13] ), .B1(n1638), 
        .C0(\matrix_b[2][13] ), .C1(n1637), .Y(n1237) );
  CLKINVX1 U1989 ( .A(n1236), .Y(n1872) );
  AOI222XL U1990 ( .A0(b33[6]), .A1(n1643), .B0(\matrix_b[6][14] ), .B1(n1638), 
        .C0(\matrix_b[2][14] ), .C1(n1637), .Y(n1236) );
  CLKINVX1 U1991 ( .A(n1235), .Y(n1873) );
  AOI222XL U1992 ( .A0(b33[7]), .A1(n1644), .B0(\matrix_b[6][15] ), .B1(n1638), 
        .C0(\matrix_b[2][15] ), .C1(n1637), .Y(n1235) );
  CLKINVX1 U1993 ( .A(n1213), .Y(n1898) );
  AOI222XL U1994 ( .A0(b32[0]), .A1(n1642), .B0(\matrix_b[6][16] ), .B1(n1640), 
        .C0(\matrix_b[1][8] ), .C1(n1206), .Y(n1213) );
  CLKINVX1 U1995 ( .A(n1212), .Y(n1899) );
  AOI222XL U1996 ( .A0(b32[1]), .A1(n1642), .B0(\matrix_b[6][17] ), .B1(n1640), 
        .C0(\matrix_b[1][9] ), .C1(n1206), .Y(n1212) );
  CLKINVX1 U1997 ( .A(n1211), .Y(n1900) );
  AOI222XL U1998 ( .A0(b32[2]), .A1(n1642), .B0(\matrix_b[6][18] ), .B1(n1640), 
        .C0(\matrix_b[1][10] ), .C1(n1206), .Y(n1211) );
  CLKINVX1 U1999 ( .A(n1210), .Y(n1901) );
  AOI222XL U2000 ( .A0(b32[3]), .A1(n1642), .B0(\matrix_b[6][19] ), .B1(n1640), 
        .C0(\matrix_b[1][11] ), .C1(n1639), .Y(n1210) );
  CLKINVX1 U2001 ( .A(n1209), .Y(n1902) );
  AOI222XL U2002 ( .A0(b32[4]), .A1(n1642), .B0(\matrix_b[6][20] ), .B1(n1640), 
        .C0(\matrix_b[1][12] ), .C1(n1639), .Y(n1209) );
  CLKINVX1 U2003 ( .A(n1208), .Y(n1903) );
  AOI222XL U2004 ( .A0(b32[5]), .A1(n1642), .B0(\matrix_b[6][21] ), .B1(n1640), 
        .C0(\matrix_b[1][13] ), .C1(n1639), .Y(n1208) );
  CLKINVX1 U2005 ( .A(n1207), .Y(n1904) );
  AOI222XL U2006 ( .A0(b32[6]), .A1(n1642), .B0(\matrix_b[6][22] ), .B1(n1640), 
        .C0(\matrix_b[1][14] ), .C1(n1639), .Y(n1207) );
  CLKINVX1 U2007 ( .A(n1204), .Y(n1905) );
  AOI222XL U2008 ( .A0(b32[7]), .A1(n1642), .B0(\matrix_b[6][23] ), .B1(n1640), 
        .C0(\matrix_b[1][15] ), .C1(n1639), .Y(n1204) );
  CLKINVX1 U2009 ( .A(n1262), .Y(n1858) );
  AOI222XL U2010 ( .A0(b24[0]), .A1(n1643), .B0(\matrix_b[5][0] ), .B1(n1638), 
        .C0(\matrix_b[3][16] ), .C1(n1637), .Y(n1262) );
  CLKINVX1 U2011 ( .A(n1261), .Y(n1859) );
  AOI222XL U2012 ( .A0(b24[1]), .A1(n1643), .B0(\matrix_b[5][1] ), .B1(n1638), 
        .C0(\matrix_b[3][17] ), .C1(n1637), .Y(n1261) );
  CLKINVX1 U2013 ( .A(n1260), .Y(n1860) );
  AOI222XL U2014 ( .A0(b24[2]), .A1(n1643), .B0(\matrix_b[5][2] ), .B1(n1215), 
        .C0(\matrix_b[3][18] ), .C1(n1637), .Y(n1260) );
  CLKINVX1 U2015 ( .A(n1259), .Y(n1861) );
  AOI222XL U2016 ( .A0(b24[3]), .A1(n1643), .B0(\matrix_b[5][3] ), .B1(n1215), 
        .C0(\matrix_b[3][19] ), .C1(n1637), .Y(n1259) );
  CLKINVX1 U2017 ( .A(n1258), .Y(n1862) );
  AOI222XL U2018 ( .A0(b24[4]), .A1(n1643), .B0(\matrix_b[5][4] ), .B1(n1215), 
        .C0(\matrix_b[3][20] ), .C1(n1637), .Y(n1258) );
  CLKINVX1 U2019 ( .A(n1257), .Y(n1863) );
  AOI222XL U2020 ( .A0(b24[5]), .A1(n1643), .B0(\matrix_b[5][5] ), .B1(n1215), 
        .C0(\matrix_b[3][21] ), .C1(n1637), .Y(n1257) );
  CLKINVX1 U2021 ( .A(n1256), .Y(n1864) );
  AOI222XL U2022 ( .A0(b24[6]), .A1(n1643), .B0(\matrix_b[5][6] ), .B1(n1638), 
        .C0(\matrix_b[3][22] ), .C1(n1637), .Y(n1256) );
  CLKINVX1 U2023 ( .A(n1255), .Y(n1865) );
  AOI222XL U2024 ( .A0(b24[7]), .A1(n1643), .B0(\matrix_b[5][7] ), .B1(n1638), 
        .C0(\matrix_b[3][23] ), .C1(n1637), .Y(n1255) );
  CLKINVX1 U2025 ( .A(n1234), .Y(n1890) );
  AOI222XL U2026 ( .A0(b23[0]), .A1(n1641), .B0(\matrix_b[5][8] ), .B1(n1640), 
        .C0(\matrix_b[2][16] ), .C1(n1639), .Y(n1234) );
  CLKINVX1 U2027 ( .A(n1233), .Y(n1891) );
  AOI222XL U2028 ( .A0(b23[1]), .A1(n1641), .B0(\matrix_b[5][9] ), .B1(n1640), 
        .C0(\matrix_b[2][17] ), .C1(n1639), .Y(n1233) );
  CLKINVX1 U2029 ( .A(n1232), .Y(n1892) );
  AOI222XL U2030 ( .A0(b23[2]), .A1(n1641), .B0(\matrix_b[5][10] ), .B1(n1205), 
        .C0(\matrix_b[2][18] ), .C1(n1639), .Y(n1232) );
  CLKINVX1 U2031 ( .A(n1231), .Y(n1893) );
  AOI222XL U2032 ( .A0(b23[3]), .A1(n1641), .B0(\matrix_b[5][11] ), .B1(n1640), 
        .C0(\matrix_b[2][19] ), .C1(n1639), .Y(n1231) );
  CLKINVX1 U2033 ( .A(n1230), .Y(n1894) );
  AOI222XL U2034 ( .A0(b23[4]), .A1(n1641), .B0(\matrix_b[5][12] ), .B1(n1640), 
        .C0(\matrix_b[2][20] ), .C1(n1639), .Y(n1230) );
  CLKINVX1 U2035 ( .A(n1229), .Y(n1895) );
  AOI222XL U2036 ( .A0(b23[5]), .A1(n1641), .B0(\matrix_b[5][13] ), .B1(n1640), 
        .C0(\matrix_b[2][21] ), .C1(n1639), .Y(n1229) );
  CLKINVX1 U2037 ( .A(n1228), .Y(n1896) );
  AOI222XL U2038 ( .A0(b23[6]), .A1(n1641), .B0(\matrix_b[5][14] ), .B1(n1640), 
        .C0(\matrix_b[2][22] ), .C1(n1206), .Y(n1228) );
  CLKINVX1 U2039 ( .A(n1227), .Y(n1897) );
  AOI222XL U2040 ( .A0(b23[7]), .A1(n1642), .B0(\matrix_b[5][15] ), .B1(n1640), 
        .C0(\matrix_b[2][23] ), .C1(n1639), .Y(n1227) );
  CLKINVX1 U2041 ( .A(n1253), .Y(n1882) );
  AOI222XL U2042 ( .A0(b14[0]), .A1(n1641), .B0(\matrix_b[4][0] ), .B1(n1205), 
        .C0(\matrix_b[3][24] ), .C1(n1639), .Y(n1253) );
  CLKINVX1 U2043 ( .A(n1252), .Y(n1883) );
  AOI222XL U2044 ( .A0(b14[1]), .A1(n1641), .B0(\matrix_b[4][1] ), .B1(n1205), 
        .C0(\matrix_b[3][25] ), .C1(n1639), .Y(n1252) );
  CLKINVX1 U2045 ( .A(n1251), .Y(n1884) );
  AOI222XL U2046 ( .A0(b14[2]), .A1(n1641), .B0(\matrix_b[4][2] ), .B1(n1205), 
        .C0(\matrix_b[3][26] ), .C1(n1639), .Y(n1251) );
  CLKINVX1 U2047 ( .A(n1250), .Y(n1885) );
  AOI222XL U2048 ( .A0(b14[3]), .A1(n1641), .B0(\matrix_b[4][3] ), .B1(n1640), 
        .C0(\matrix_b[3][27] ), .C1(n1639), .Y(n1250) );
  CLKINVX1 U2049 ( .A(n1249), .Y(n1886) );
  AOI222XL U2050 ( .A0(b14[4]), .A1(n1641), .B0(\matrix_b[4][4] ), .B1(n1640), 
        .C0(\matrix_b[3][28] ), .C1(n1639), .Y(n1249) );
  CLKINVX1 U2051 ( .A(n1248), .Y(n1887) );
  AOI222XL U2052 ( .A0(b14[5]), .A1(n1641), .B0(\matrix_b[4][5] ), .B1(n1640), 
        .C0(\matrix_b[3][29] ), .C1(n1639), .Y(n1248) );
  CLKINVX1 U2053 ( .A(n1247), .Y(n1888) );
  AOI222XL U2054 ( .A0(b14[6]), .A1(n1641), .B0(\matrix_b[4][6] ), .B1(n1640), 
        .C0(\matrix_b[3][30] ), .C1(n1639), .Y(n1247) );
  CLKINVX1 U2055 ( .A(n1246), .Y(n1889) );
  AOI222XL U2056 ( .A0(b14[7]), .A1(n1641), .B0(\matrix_b[4][7] ), .B1(n1640), 
        .C0(\matrix_b[3][31] ), .C1(n1639), .Y(n1246) );
  CLKINVX1 U2057 ( .A(n1223), .Y(n1874) );
  AOI222XL U2058 ( .A0(b42[0]), .A1(n1644), .B0(\matrix_b[7][16] ), .B1(n1638), 
        .C0(\matrix_b[1][0] ), .C1(n1216), .Y(n1223) );
  CLKINVX1 U2059 ( .A(n1222), .Y(n1875) );
  AOI222XL U2060 ( .A0(b42[1]), .A1(n1644), .B0(\matrix_b[7][17] ), .B1(n1638), 
        .C0(\matrix_b[1][1] ), .C1(n1216), .Y(n1222) );
  CLKINVX1 U2061 ( .A(n1221), .Y(n1876) );
  AOI222XL U2062 ( .A0(b42[2]), .A1(n1644), .B0(\matrix_b[7][18] ), .B1(n1638), 
        .C0(\matrix_b[1][2] ), .C1(n1216), .Y(n1221) );
  CLKINVX1 U2063 ( .A(n1220), .Y(n1877) );
  AOI222XL U2064 ( .A0(b42[3]), .A1(n1644), .B0(\matrix_b[7][19] ), .B1(n1638), 
        .C0(\matrix_b[1][3] ), .C1(n1216), .Y(n1220) );
  CLKINVX1 U2065 ( .A(n1219), .Y(n1878) );
  AOI222XL U2066 ( .A0(b42[4]), .A1(n1644), .B0(\matrix_b[7][20] ), .B1(n1638), 
        .C0(\matrix_b[1][4] ), .C1(n1637), .Y(n1219) );
  CLKINVX1 U2067 ( .A(n1218), .Y(n1879) );
  AOI222XL U2068 ( .A0(b42[5]), .A1(n1644), .B0(\matrix_b[7][21] ), .B1(n1638), 
        .C0(\matrix_b[1][5] ), .C1(n1637), .Y(n1218) );
  CLKINVX1 U2069 ( .A(n1217), .Y(n1880) );
  AOI222XL U2070 ( .A0(b42[6]), .A1(n1644), .B0(\matrix_b[7][22] ), .B1(n1638), 
        .C0(\matrix_b[1][6] ), .C1(n1637), .Y(n1217) );
  CLKINVX1 U2071 ( .A(n1214), .Y(n1881) );
  AOI222XL U2072 ( .A0(b42[7]), .A1(n1644), .B0(\matrix_b[7][23] ), .B1(n1638), 
        .C0(\matrix_b[1][7] ), .C1(n1637), .Y(n1214) );
  CLKINVX1 U2073 ( .A(w24[0]), .Y(n1786) );
  CLKINVX1 U2074 ( .A(w34[0]), .Y(n1794) );
  CLKINVX1 U2075 ( .A(w14[0]), .Y(n1770) );
  CLKINVX1 U2076 ( .A(w24[1]), .Y(n1785) );
  CLKINVX1 U2077 ( .A(w24[2]), .Y(n1784) );
  CLKINVX1 U2078 ( .A(w24[3]), .Y(n1783) );
  CLKINVX1 U2079 ( .A(w34[1]), .Y(n1793) );
  CLKINVX1 U2080 ( .A(w34[2]), .Y(n1792) );
  CLKINVX1 U2081 ( .A(w34[3]), .Y(n1791) );
  CLKINVX1 U2082 ( .A(w14[1]), .Y(n1769) );
  CLKINVX1 U2083 ( .A(w14[2]), .Y(n1768) );
  CLKINVX1 U2084 ( .A(w14[3]), .Y(n1767) );
  CLKBUFX3 U2085 ( .A(index_a[3]), .Y(n1694) );
  CLKBUFX3 U2086 ( .A(index_b[3]), .Y(n1687) );
  CLKBUFX3 U2087 ( .A(n964), .Y(n1669) );
  NAND3X1 U2088 ( .A(n1629), .B(n700), .C(n1164), .Y(n964) );
  NAND3X1 U2089 ( .A(n1628), .B(n699), .C(n1197), .Y(n972) );
  NAND3X1 U2090 ( .A(n1628), .B(n699), .C(n1165), .Y(n968) );
  CLKBUFX3 U2091 ( .A(index_a[4]), .Y(n1695) );
  CLKBUFX3 U2092 ( .A(index_b[4]), .Y(n1688) );
  NAND4X1 U2093 ( .A(l[2]), .B(n957), .C(n631), .D(n630), .Y(n843) );
  NOR2X1 U2094 ( .A(cur_state[0]), .B(cur_state[1]), .Y(n1509) );
  CLKINVX1 U2095 ( .A(w44[4]), .Y(n1798) );
  CLKINVX1 U2096 ( .A(w44[5]), .Y(n1797) );
  CLKINVX1 U2097 ( .A(w44[6]), .Y(n1796) );
  CLKINVX1 U2098 ( .A(w44[7]), .Y(n1795) );
  CLKINVX1 U2099 ( .A(w24[4]), .Y(n1782) );
  CLKINVX1 U2100 ( .A(w24[5]), .Y(n1781) );
  CLKINVX1 U2101 ( .A(w24[6]), .Y(n1780) );
  CLKINVX1 U2102 ( .A(w24[7]), .Y(n1779) );
  CLKINVX1 U2103 ( .A(w34[4]), .Y(n1790) );
  CLKINVX1 U2104 ( .A(w34[5]), .Y(n1789) );
  CLKINVX1 U2105 ( .A(w34[6]), .Y(n1788) );
  CLKINVX1 U2106 ( .A(w34[7]), .Y(n1787) );
  CLKINVX1 U2107 ( .A(w14[4]), .Y(n1766) );
  CLKINVX1 U2108 ( .A(w14[5]), .Y(n1765) );
  CLKINVX1 U2109 ( .A(w14[6]), .Y(n1764) );
  CLKINVX1 U2110 ( .A(w14[7]), .Y(n1763) );
  OAI2BB1X1 U2111 ( .A0N(cur_state[0]), .A1N(load_en), .B0(n163), .Y(
        next_state[1]) );
  CLKBUFX3 U2112 ( .A(data_out_a[8]), .Y(n1578) );
  CLKBUFX3 U2113 ( .A(data_out_a[9]), .Y(n1579) );
  CLKBUFX3 U2114 ( .A(data_out_a[10]), .Y(n1580) );
  CLKBUFX3 U2115 ( .A(data_out_a[11]), .Y(n1581) );
  CLKBUFX3 U2116 ( .A(data_out_a[12]), .Y(n1582) );
  CLKBUFX3 U2117 ( .A(data_out_a[13]), .Y(n1583) );
  CLKBUFX3 U2118 ( .A(data_out_a[14]), .Y(n1584) );
  CLKBUFX3 U2119 ( .A(data_out_a[15]), .Y(n1585) );
  CLKBUFX3 U2120 ( .A(data_out_a[16]), .Y(n1586) );
  CLKBUFX3 U2121 ( .A(data_out_a[17]), .Y(n1587) );
  CLKBUFX3 U2122 ( .A(data_out_a[18]), .Y(n1588) );
  CLKBUFX3 U2123 ( .A(data_out_a[19]), .Y(n1589) );
  CLKBUFX3 U2124 ( .A(data_out_a[20]), .Y(n1590) );
  CLKBUFX3 U2125 ( .A(data_out_a[21]), .Y(n1591) );
  CLKBUFX3 U2126 ( .A(data_out_a[22]), .Y(n1592) );
  CLKBUFX3 U2127 ( .A(data_out_a[23]), .Y(n1593) );
  CLKINVX1 U2128 ( .A(n1521), .Y(n1851) );
  NOR4X1 U2129 ( .A(n1626), .B(n1627), .C(n1628), .D(n1621), .Y(n1697) );
  NOR4X1 U2130 ( .A(n1622), .B(n1623), .C(n1624), .D(n1625), .Y(n1696) );
  NOR3X1 U2131 ( .A(n1624), .B(n1622), .C(n1623), .Y(n1700) );
  AND3X1 U2132 ( .A(n1630), .B(n1631), .C(n1629), .Y(n1698) );
  NOR4X1 U2133 ( .A(n1627), .B(n1628), .C(n1621), .D(n1698), .Y(n1699) );
  OR2X1 U2134 ( .A(n1622), .B(n1623), .Y(n1701) );
  OR4X1 U2135 ( .A(n1625), .B(n1626), .C(n1624), .D(n1701), .Y(n1703) );
  AO21X1 U2136 ( .A0(n1629), .A1(n1630), .B0(n1621), .Y(n1702) );
  NOR3X1 U2137 ( .A(n1624), .B(n1622), .C(n1623), .Y(n1706) );
  OA21XL U2138 ( .A0(n1630), .A1(n1631), .B0(n1629), .Y(n1704) );
  NOR4X1 U2139 ( .A(n1627), .B(n1621), .C(n1628), .D(n1704), .Y(n1705) );
  NOR2BX1 U2140 ( .AN(N783), .B(n1627), .Y(n1714) );
  NAND2BX1 U2141 ( .AN(N781), .B(n1629), .Y(n1709) );
  OAI21XL U2142 ( .A0(N780), .A1(n1743), .B0(n1707), .Y(n1712) );
  NOR2BX1 U2143 ( .AN(N781), .B(n1629), .Y(n1708) );
  OR4X1 U2144 ( .A(n1624), .B(n1625), .C(n1622), .D(n1623), .Y(n1715) );
  NOR2BX1 U2145 ( .AN(N715), .B(n1627), .Y(n1725) );
  NAND2BX1 U2146 ( .AN(N713), .B(n1629), .Y(n1720) );
  OAI21XL U2147 ( .A0(N712), .A1(n1743), .B0(n1718), .Y(n1723) );
  NOR2BX1 U2148 ( .AN(N713), .B(n1629), .Y(n1719) );
  OAI22XL U2149 ( .A0(n1725), .A1(n1724), .B0(N715), .B1(n1533), .Y(n1727) );
  OR4X1 U2150 ( .A(n1624), .B(n1625), .C(n1622), .D(n1623), .Y(n1726) );
  NAND2X1 U2151 ( .A(n1629), .B(n1744), .Y(n1730) );
  NOR2BX1 U2152 ( .AN(n1626), .B(n1573), .Y(n1729) );
  NOR4X1 U2153 ( .A(n1625), .B(n1729), .C(n1623), .D(n1624), .Y(n1738) );
  OAI21XL U2154 ( .A0(N789), .A1(n1533), .B0(n1738), .Y(n1741) );
  NOR2X1 U2155 ( .A(n1529), .B(n1631), .Y(n1732) );
  OAI211X1 U2156 ( .A0(N789), .A1(n1533), .B0(n1735), .C0(n1734), .Y(n1736) );
  OAI221XL U2157 ( .A0(n1627), .A1(n1746), .B0(n1626), .B1(n1747), .C0(n1736), 
        .Y(n1737) );
  AND4X1 U2158 ( .A(n1738), .B(n1737), .C(n1516), .D(n1519), .Y(N791) );
  NAND2X1 U2159 ( .A(n1631), .B(n1529), .Y(n1739) );
  AOI22X1 U2160 ( .A0(n1739), .A1(n1743), .B0(n1739), .B1(N786), .Y(n1740) );
  NOR4X1 U2161 ( .A(n1742), .B(n1741), .C(N791), .D(n1740), .Y(N793) );
endmodule

